--
-- DVB IP
--
-- Copyright 2020 by Suoto <andre820@gmail.com>
--
-- This file is part of the DVB IP.
--
-- DVB IP is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- DVB IP is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with DVB IP.  If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library fpga_cores;
use fpga_cores.common_pkg.all;

use work.dvb_utils_pkg.all;

-- Summary of statistics

--    table                               depth    width (bits)    width (entries)    total (bytes)    18k BRAMs    36k BRAMs
----  --------------------------------  -------  --------------  -----------------  ---------------  -----------  -----------
--    ldpc_table_FECFRAME_NORMAL_C1_2        90             115                  9             1294            7            4
--    ldpc_table_FECFRAME_NORMAL_C1_3        60             196                 13             1470           11            6
--    ldpc_table_FECFRAME_NORMAL_C1_4        45             196                 13             1103           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_3       120             189                 14             2835           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_5        72             196                 13             1764           11            6
--    ldpc_table_FECFRAME_NORMAL_C3_4       135             164                 13             2768           10            5
--    ldpc_table_FECFRAME_NORMAL_C3_5       108             184                 13             2484           11            6
--    ldpc_table_FECFRAME_NORMAL_C4_5       144             150                 12             2700            9            5
--    ldpc_table_FECFRAME_NORMAL_C5_6       150             177                 14             3319           10            5
--    ldpc_table_FECFRAME_NORMAL_C8_9       160              46                  5              920            3            2
--    ldpc_table_FECFRAME_NORMAL_C9_10      162              46                  5              932            3            2
--    ldpc_table_FECFRAME_SHORT_C1_2         20             100                  9              250            6            3
--    ldpc_table_FECFRAME_SHORT_C1_3         15             170                 13              319           10            5
--    ldpc_table_FECFRAME_SHORT_C1_4          9             171                 13              193           10            5
--    ldpc_table_FECFRAME_SHORT_C2_3         30             156                 14              585            9            5
--    ldpc_table_FECFRAME_SHORT_C2_5         18             168                 13              378           10            5
--    ldpc_table_FECFRAME_SHORT_C3_4         33             133                 13              549            8            4
--    ldpc_table_FECFRAME_SHORT_C3_5         27             160                 13              540            9            5
--    ldpc_table_FECFRAME_SHORT_C4_5         35              30                  4              132            2            1
--    ldpc_table_FECFRAME_SHORT_C5_6         37             139                 14              643            8            4
--    ldpc_table_FECFRAME_SHORT_C8_9         40              37                  5              185            3            2

package ldpc_tables_pkg is


  -- LDPC_TABLE_FECFRAME_<frame_length>_<code_rate>_COLUMN_WIDTHS constants have the bit
  -- width of each row

  -- LDPC_TABLE_FECFRAME_<frame_length>_<code_rate> is the actual LDPC where the number of
  -- columns is normalized to the row with most columns and the first column of each row
  -- contains the number of valid elements within the row. Elements outisde the valid range
  -- are represented as -1


  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_2.csv, table is 90x115 (1293.75 bytes)
  -- Resource estimation: 7 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 7, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2 : integer_2d_array_t(0 to 89)(0 to 8) := (
    0 => integer_vector_t'(0 => 8, 1 => 54, 2 => 9318, 3 => 14392, 4 => 27561, 5 => 26909, 6 => 10219, 7 => 2534, 8 => 8597),
    1 => integer_vector_t'(0 => 8, 1 => 55, 2 => 7263, 3 => 4635, 4 => 2530, 5 => 28130, 6 => 3033, 7 => 23830, 8 => 3651),
    2 => integer_vector_t'(0 => 8, 1 => 56, 2 => 24731, 3 => 23583, 4 => 26036, 5 => 17299, 6 => 5750, 7 => 792, 8 => 9169),
    3 => integer_vector_t'(0 => 8, 1 => 57, 2 => 5811, 3 => 26154, 4 => 18653, 5 => 11551, 6 => 15447, 7 => 13685, 8 => 16264),
    4 => integer_vector_t'(0 => 8, 1 => 58, 2 => 12610, 3 => 11347, 4 => 28768, 5 => 2792, 6 => 3174, 7 => 29371, 8 => 12997),
    5 => integer_vector_t'(0 => 8, 1 => 59, 2 => 16789, 3 => 16018, 4 => 21449, 5 => 6165, 6 => 21202, 7 => 15850, 8 => 3186),
    6 => integer_vector_t'(0 => 8, 1 => 60, 2 => 31016, 3 => 21449, 4 => 17618, 5 => 6213, 6 => 12166, 7 => 8334, 8 => 18212),
    7 => integer_vector_t'(0 => 8, 1 => 61, 2 => 22836, 3 => 14213, 4 => 11327, 5 => 5896, 6 => 718, 7 => 11727, 8 => 9308),
    8 => integer_vector_t'(0 => 8, 1 => 62, 2 => 2091, 3 => 24941, 4 => 29966, 5 => 23634, 6 => 9013, 7 => 15587, 8 => 5444),
    9 => integer_vector_t'(0 => 8, 1 => 63, 2 => 22207, 3 => 3983, 4 => 16904, 5 => 28534, 6 => 21415, 7 => 27524, 8 => 25912),
    10 => integer_vector_t'(0 => 8, 1 => 64, 2 => 25687, 3 => 4501, 4 => 22193, 5 => 14665, 6 => 14798, 7 => 16158, 8 => 5491),
    11 => integer_vector_t'(0 => 8, 1 => 65, 2 => 4520, 3 => 17094, 4 => 23397, 5 => 4264, 6 => 22370, 7 => 16941, 8 => 21526),
    12 => integer_vector_t'(0 => 8, 1 => 66, 2 => 10490, 3 => 6182, 4 => 32370, 5 => 9597, 6 => 30841, 7 => 25954, 8 => 2762),
    13 => integer_vector_t'(0 => 8, 1 => 67, 2 => 22120, 3 => 22865, 4 => 29870, 5 => 15147, 6 => 13668, 7 => 14955, 8 => 19235),
    14 => integer_vector_t'(0 => 8, 1 => 68, 2 => 6689, 3 => 18408, 4 => 18346, 5 => 9918, 6 => 25746, 7 => 5443, 8 => 20645),
    15 => integer_vector_t'(0 => 8, 1 => 69, 2 => 29982, 3 => 12529, 4 => 13858, 5 => 4746, 6 => 30370, 7 => 10023, 8 => 24828),
    16 => integer_vector_t'(0 => 8, 1 => 70, 2 => 1262, 3 => 28032, 4 => 29888, 5 => 13063, 6 => 24033, 7 => 21951, 8 => 7863),
    17 => integer_vector_t'(0 => 8, 1 => 71, 2 => 6594, 3 => 29642, 4 => 31451, 5 => 14831, 6 => 9509, 7 => 9335, 8 => 31552),
    18 => integer_vector_t'(0 => 8, 1 => 72, 2 => 1358, 3 => 6454, 4 => 16633, 5 => 20354, 6 => 24598, 7 => 624, 8 => 5265),
    19 => integer_vector_t'(0 => 8, 1 => 73, 2 => 19529, 3 => 295, 4 => 18011, 5 => 3080, 6 => 13364, 7 => 8032, 8 => 15323),
    20 => integer_vector_t'(0 => 8, 1 => 74, 2 => 11981, 3 => 1510, 4 => 7960, 5 => 21462, 6 => 9129, 7 => 11370, 8 => 25741),
    21 => integer_vector_t'(0 => 8, 1 => 75, 2 => 9276, 3 => 29656, 4 => 4543, 5 => 30699, 6 => 20646, 7 => 21921, 8 => 28050),
    22 => integer_vector_t'(0 => 8, 1 => 76, 2 => 15975, 3 => 25634, 4 => 5520, 5 => 31119, 6 => 13715, 7 => 21949, 8 => 19605),
    23 => integer_vector_t'(0 => 8, 1 => 77, 2 => 18688, 3 => 4608, 4 => 31755, 5 => 30165, 6 => 13103, 7 => 10706, 8 => 29224),
    24 => integer_vector_t'(0 => 8, 1 => 78, 2 => 21514, 3 => 23117, 4 => 12245, 5 => 26035, 6 => 31656, 7 => 25631, 8 => 30699),
    25 => integer_vector_t'(0 => 8, 1 => 79, 2 => 9674, 3 => 24966, 4 => 31285, 5 => 29908, 6 => 17042, 7 => 24588, 8 => 31857),
    26 => integer_vector_t'(0 => 8, 1 => 80, 2 => 21856, 3 => 27777, 4 => 29919, 5 => 27000, 6 => 14897, 7 => 11409, 8 => 7122),
    27 => integer_vector_t'(0 => 8, 1 => 81, 2 => 29773, 3 => 23310, 4 => 263, 5 => 4877, 6 => 28622, 7 => 20545, 8 => 22092),
    28 => integer_vector_t'(0 => 8, 1 => 82, 2 => 15605, 3 => 5651, 4 => 21864, 5 => 3967, 6 => 14419, 7 => 22757, 8 => 15896),
    29 => integer_vector_t'(0 => 8, 1 => 83, 2 => 30145, 3 => 1759, 4 => 10139, 5 => 29223, 6 => 26086, 7 => 10556, 8 => 5098),
    30 => integer_vector_t'(0 => 8, 1 => 84, 2 => 18815, 3 => 16575, 4 => 2936, 5 => 24457, 6 => 26738, 7 => 6030, 8 => 505),
    31 => integer_vector_t'(0 => 8, 1 => 85, 2 => 30326, 3 => 22298, 4 => 27562, 5 => 20131, 6 => 26390, 7 => 6247, 8 => 24791),
    32 => integer_vector_t'(0 => 8, 1 => 86, 2 => 928, 3 => 29246, 4 => 21246, 5 => 12400, 6 => 15311, 7 => 32309, 8 => 18608),
    33 => integer_vector_t'(0 => 8, 1 => 87, 2 => 20314, 3 => 6025, 4 => 26689, 5 => 16302, 6 => 2296, 7 => 3244, 8 => 19613),
    34 => integer_vector_t'(0 => 8, 1 => 88, 2 => 6237, 3 => 11943, 4 => 22851, 5 => 15642, 6 => 23857, 7 => 15112, 8 => 20947),
    35 => integer_vector_t'(0 => 8, 1 => 89, 2 => 26403, 3 => 25168, 4 => 19038, 5 => 18384, 6 => 8882, 7 => 12719, 8 => 7093),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 14567, 3 => 24965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3908, 3 => 100, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10279, 3 => 240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 24102, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 12383, 3 => 4173, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 13861, 3 => 15918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 21327, 3 => 1046, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5288, 3 => 14579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 28158, 3 => 8069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 16583, 3 => 11098, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 16681, 3 => 28363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 13980, 3 => 24725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 32169, 3 => 17989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 10907, 3 => 2767, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 21557, 3 => 3818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 26676, 3 => 12422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 7676, 3 => 8754, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 14905, 3 => 20232, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 15719, 3 => 24646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 31942, 3 => 8589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 19978, 3 => 27197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 27060, 3 => 15071, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6071, 3 => 26649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10393, 3 => 11176, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 9597, 3 => 13370, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7081, 3 => 17677, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 1433, 3 => 19513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 26925, 3 => 9014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 19202, 3 => 8900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 18152, 3 => 30647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20803, 3 => 1737, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 11804, 3 => 25221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 31683, 3 => 17783, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 29694, 3 => 9345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 12280, 3 => 26611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 6526, 3 => 26122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 26165, 3 => 11241, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 7666, 3 => 26962, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 16290, 3 => 8480, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 11774, 3 => 10120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 30051, 3 => 30426, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 1335, 3 => 15424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6865, 3 => 17742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 31779, 3 => 12489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 32120, 3 => 21001, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 14508, 3 => 6996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 979, 3 => 25024, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 4554, 3 => 21896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 7989, 3 => 21777, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 4972, 3 => 20661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 6612, 3 => 2730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 12742, 3 => 4418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 29194, 3 => 595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 19267, 3 => 20113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_3.csv, table is 60x196 (1470.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3 : integer_2d_array_t(0 to 59)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 34903, 2 => 20927, 3 => 32093, 4 => 1052, 5 => 25611, 6 => 16093, 7 => 16454, 8 => 5520, 9 => 506, 10 => 37399, 11 => 18518, 12 => 21120),
    1 => integer_vector_t'(0 => 12, 1 => 11636, 2 => 14594, 3 => 22158, 4 => 14763, 5 => 15333, 6 => 6838, 7 => 22222, 8 => 37856, 9 => 14985, 10 => 31041, 11 => 18704, 12 => 32910),
    2 => integer_vector_t'(0 => 12, 1 => 17449, 2 => 1665, 3 => 35639, 4 => 16624, 5 => 12867, 6 => 12449, 7 => 10241, 8 => 11650, 9 => 25622, 10 => 34372, 11 => 19878, 12 => 26894),
    3 => integer_vector_t'(0 => 12, 1 => 29235, 2 => 19780, 3 => 36056, 4 => 20129, 5 => 20029, 6 => 5457, 7 => 8157, 8 => 35554, 9 => 21237, 10 => 7943, 11 => 13873, 12 => 14980),
    4 => integer_vector_t'(0 => 12, 1 => 9912, 2 => 7143, 3 => 35911, 4 => 12043, 5 => 17360, 6 => 37253, 7 => 25588, 8 => 11827, 9 => 29152, 10 => 21936, 11 => 24125, 12 => 40870),
    5 => integer_vector_t'(0 => 12, 1 => 40701, 2 => 36035, 3 => 39556, 4 => 12366, 5 => 19946, 6 => 29072, 7 => 16365, 8 => 35495, 9 => 22686, 10 => 11106, 11 => 8756, 12 => 34863),
    6 => integer_vector_t'(0 => 12, 1 => 19165, 2 => 15702, 3 => 13536, 4 => 40238, 5 => 4465, 6 => 40034, 7 => 40590, 8 => 37540, 9 => 17162, 10 => 1712, 11 => 20577, 12 => 14138),
    7 => integer_vector_t'(0 => 12, 1 => 31338, 2 => 19342, 3 => 9301, 4 => 39375, 5 => 3211, 6 => 1316, 7 => 33409, 8 => 28670, 9 => 12282, 10 => 6118, 11 => 29236, 12 => 35787),
    8 => integer_vector_t'(0 => 12, 1 => 11504, 2 => 30506, 3 => 19558, 4 => 5100, 5 => 24188, 6 => 24738, 7 => 30397, 8 => 33775, 9 => 9699, 10 => 6215, 11 => 3397, 12 => 37451),
    9 => integer_vector_t'(0 => 12, 1 => 34689, 2 => 23126, 3 => 7571, 4 => 1058, 5 => 12127, 6 => 27518, 7 => 23064, 8 => 11265, 9 => 14867, 10 => 30451, 11 => 28289, 12 => 2966),
    10 => integer_vector_t'(0 => 12, 1 => 11660, 2 => 15334, 3 => 16867, 4 => 15160, 5 => 38343, 6 => 3778, 7 => 4265, 8 => 39139, 9 => 17293, 10 => 26229, 11 => 42604, 12 => 13486),
    11 => integer_vector_t'(0 => 12, 1 => 31497, 2 => 1365, 3 => 14828, 4 => 7453, 5 => 26350, 6 => 41346, 7 => 28643, 8 => 23421, 9 => 8354, 10 => 16255, 11 => 11055, 12 => 24279),
    12 => integer_vector_t'(0 => 12, 1 => 15687, 2 => 12467, 3 => 13906, 4 => 5215, 5 => 41328, 6 => 23755, 7 => 20800, 8 => 6447, 9 => 7970, 10 => 2803, 11 => 33262, 12 => 39843),
    13 => integer_vector_t'(0 => 12, 1 => 5363, 2 => 22469, 3 => 38091, 4 => 28457, 5 => 36696, 6 => 34471, 7 => 23619, 8 => 2404, 9 => 24229, 10 => 41754, 11 => 1297, 12 => 18563),
    14 => integer_vector_t'(0 => 12, 1 => 3673, 2 => 39070, 3 => 14480, 4 => 30279, 5 => 37483, 6 => 7580, 7 => 29519, 8 => 30519, 9 => 39831, 10 => 20252, 11 => 18132, 12 => 20010),
    15 => integer_vector_t'(0 => 12, 1 => 34386, 2 => 7252, 3 => 27526, 4 => 12950, 5 => 6875, 6 => 43020, 7 => 31566, 8 => 39069, 9 => 18985, 10 => 15541, 11 => 40020, 12 => 16715),
    16 => integer_vector_t'(0 => 12, 1 => 1721, 2 => 37332, 3 => 39953, 4 => 17430, 5 => 32134, 6 => 29162, 7 => 10490, 8 => 12971, 9 => 28581, 10 => 29331, 11 => 6489, 12 => 35383),
    17 => integer_vector_t'(0 => 12, 1 => 736, 2 => 7022, 3 => 42349, 4 => 8783, 5 => 6767, 6 => 11871, 7 => 21675, 8 => 10325, 9 => 11548, 10 => 25978, 11 => 431, 12 => 24085),
    18 => integer_vector_t'(0 => 12, 1 => 1925, 2 => 10602, 3 => 28585, 4 => 12170, 5 => 15156, 6 => 34404, 7 => 8351, 8 => 13273, 9 => 20208, 10 => 5800, 11 => 15367, 12 => 21764),
    19 => integer_vector_t'(0 => 12, 1 => 16279, 2 => 37832, 3 => 34792, 4 => 21250, 5 => 34192, 6 => 7406, 7 => 41488, 8 => 18346, 9 => 29227, 10 => 26127, 11 => 25493, 12 => 7048),
    20 => integer_vector_t'(0 => 3, 1 => 39948, 2 => 28229, 3 => 24899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 17408, 2 => 14274, 3 => 38993, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 38774, 2 => 15968, 3 => 28459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 41404, 2 => 27249, 3 => 27425, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 41229, 2 => 6082, 3 => 43114, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 13957, 2 => 4979, 3 => 40654, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 3093, 2 => 3438, 3 => 34992, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 34082, 2 => 6172, 3 => 28760, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 42210, 2 => 34141, 3 => 41021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14705, 2 => 17783, 3 => 10134, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 41755, 2 => 39884, 3 => 22773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14615, 2 => 15593, 3 => 1642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 29111, 2 => 37061, 3 => 39860, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 9579, 2 => 33552, 3 => 633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 12951, 2 => 21137, 3 => 39608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 38244, 2 => 27361, 3 => 29417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 2939, 2 => 10172, 3 => 36479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 29094, 2 => 5357, 3 => 19224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 9562, 2 => 24436, 3 => 28637, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 40177, 2 => 2326, 3 => 13504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 6834, 2 => 21583, 3 => 42516, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 40651, 2 => 42810, 3 => 25709, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 31557, 2 => 32138, 3 => 38142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 18624, 2 => 41867, 3 => 39296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 37560, 2 => 14295, 3 => 16245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 6821, 2 => 21679, 3 => 31570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 25339, 2 => 25083, 3 => 22081, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 8047, 2 => 697, 3 => 35268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 9884, 2 => 17073, 3 => 19995, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 26848, 2 => 35245, 3 => 8390, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 18658, 2 => 16134, 3 => 14807, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 12201, 2 => 32944, 3 => 5035, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 25236, 2 => 1216, 3 => 38986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 42994, 2 => 24782, 3 => 8681, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 28321, 2 => 4932, 3 => 34249, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 4107, 2 => 29382, 3 => 32124, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 22157, 2 => 2624, 3 => 14468, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 38788, 2 => 27081, 3 => 7936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4368, 2 => 26148, 3 => 10578, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 25353, 2 => 4122, 3 => 39751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_4.csv, table is 45x196 (1102.5 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4 : integer_2d_array_t(0 to 44)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 23606, 2 => 36098, 3 => 1140, 4 => 28859, 5 => 18148, 6 => 18510, 7 => 6226, 8 => 540, 9 => 42014, 10 => 20879, 11 => 23802, 12 => 47088),
    1 => integer_vector_t'(0 => 12, 1 => 16419, 2 => 24928, 3 => 16609, 4 => 17248, 5 => 7693, 6 => 24997, 7 => 42587, 8 => 16858, 9 => 34921, 10 => 21042, 11 => 37024, 12 => 20692),
    2 => integer_vector_t'(0 => 12, 1 => 1874, 2 => 40094, 3 => 18704, 4 => 14474, 5 => 14004, 6 => 11519, 7 => 13106, 8 => 28826, 9 => 38669, 10 => 22363, 11 => 30255, 12 => 31105),
    3 => integer_vector_t'(0 => 12, 1 => 22254, 2 => 40564, 3 => 22645, 4 => 22532, 5 => 6134, 6 => 9176, 7 => 39998, 8 => 23892, 9 => 8937, 10 => 15608, 11 => 16854, 12 => 31009),
    4 => integer_vector_t'(0 => 12, 1 => 8037, 2 => 40401, 3 => 13550, 4 => 19526, 5 => 41902, 6 => 28782, 7 => 13304, 8 => 32796, 9 => 24679, 10 => 27140, 11 => 45980, 12 => 10021),
    5 => integer_vector_t'(0 => 12, 1 => 40540, 2 => 44498, 3 => 13911, 4 => 22435, 5 => 32701, 6 => 18405, 7 => 39929, 8 => 25521, 9 => 12497, 10 => 9851, 11 => 39223, 12 => 34823),
    6 => integer_vector_t'(0 => 12, 1 => 15233, 2 => 45333, 3 => 5041, 4 => 44979, 5 => 45710, 6 => 42150, 7 => 19416, 8 => 1892, 9 => 23121, 10 => 15860, 11 => 8832, 12 => 10308),
    7 => integer_vector_t'(0 => 12, 1 => 10468, 2 => 44296, 3 => 3611, 4 => 1480, 5 => 37581, 6 => 32254, 7 => 13817, 8 => 6883, 9 => 32892, 10 => 40258, 11 => 46538, 12 => 11940),
    8 => integer_vector_t'(0 => 12, 1 => 6705, 2 => 21634, 3 => 28150, 4 => 43757, 5 => 895, 6 => 6547, 7 => 20970, 8 => 28914, 9 => 30117, 10 => 25736, 11 => 41734, 12 => 11392),
    9 => integer_vector_t'(0 => 12, 1 => 22002, 2 => 5739, 3 => 27210, 4 => 27828, 5 => 34192, 6 => 37992, 7 => 10915, 8 => 6998, 9 => 3824, 10 => 42130, 11 => 4494, 12 => 35739),
    10 => integer_vector_t'(0 => 12, 1 => 8515, 2 => 1191, 3 => 13642, 4 => 30950, 5 => 25943, 6 => 12673, 7 => 16726, 8 => 34261, 9 => 31828, 10 => 3340, 11 => 8747, 12 => 39225),
    11 => integer_vector_t'(0 => 12, 1 => 18979, 2 => 17058, 3 => 43130, 4 => 4246, 5 => 4793, 6 => 44030, 7 => 19454, 8 => 29511, 9 => 47929, 10 => 15174, 11 => 24333, 12 => 19354),
    12 => integer_vector_t'(0 => 12, 1 => 16694, 2 => 8381, 3 => 29642, 4 => 46516, 5 => 32224, 6 => 26344, 7 => 9405, 8 => 18292, 9 => 12437, 10 => 27316, 11 => 35466, 12 => 41992),
    13 => integer_vector_t'(0 => 12, 1 => 15642, 2 => 5871, 3 => 46489, 4 => 26723, 5 => 23396, 6 => 7257, 7 => 8974, 8 => 3156, 9 => 37420, 10 => 44823, 11 => 35423, 12 => 13541),
    14 => integer_vector_t'(0 => 12, 1 => 42858, 2 => 32008, 3 => 41282, 4 => 38773, 5 => 26570, 6 => 2702, 7 => 27260, 8 => 46974, 9 => 1469, 10 => 20887, 11 => 27426, 12 => 38553),
    15 => integer_vector_t'(0 => 3, 1 => 22152, 2 => 24261, 3 => 8297, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 19347, 2 => 9978, 3 => 27802, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 34991, 2 => 6354, 3 => 33561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 29782, 2 => 30875, 3 => 29523, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 9278, 2 => 48512, 3 => 14349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 38061, 2 => 4165, 3 => 43878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 8548, 2 => 33172, 3 => 34410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22535, 2 => 28811, 3 => 23950, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 20439, 2 => 4027, 3 => 24186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 38618, 2 => 8187, 3 => 30947, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 35538, 2 => 43880, 3 => 21459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 7091, 2 => 45616, 3 => 15063, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 5505, 2 => 9315, 3 => 21908, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 36046, 2 => 32914, 3 => 11836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 7304, 2 => 39782, 3 => 33721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 16905, 2 => 29962, 3 => 12980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11171, 2 => 23709, 3 => 22460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 34541, 2 => 9937, 3 => 44500, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 14035, 2 => 47316, 3 => 8815, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 15057, 2 => 45482, 3 => 24461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 30518, 2 => 36877, 3 => 879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7583, 2 => 13364, 3 => 24332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 448, 2 => 27056, 3 => 4682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 12083, 2 => 31378, 3 => 21670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 1159, 2 => 18031, 3 => 2221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 17028, 2 => 38715, 3 => 9350, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 17343, 2 => 24530, 3 => 29574, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 46128, 2 => 31039, 3 => 32818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 20373, 2 => 36967, 3 => 18345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 46685, 2 => 20622, 3 => 32806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_3.csv, table is 120x189 (2835.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 14, 9 => 15, 10 => 15, 11 => 15, 12 => 15, 13 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3 : integer_2d_array_t(0 to 119)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 10491, 3 => 16043, 4 => 506, 5 => 12826, 6 => 8065, 7 => 8226, 8 => 2767, 9 => 240, 10 => 18673, 11 => 9279, 12 => 10579, 13 => 20928),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 17819, 3 => 8313, 4 => 6433, 5 => 6224, 6 => 5120, 7 => 5824, 8 => 12812, 9 => 17187, 10 => 9940, 11 => 13447, 12 => 13825, 13 => 18483),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 17957, 3 => 6024, 4 => 8681, 5 => 18628, 6 => 12794, 7 => 5915, 8 => 14576, 9 => 10970, 10 => 12064, 11 => 20437, 12 => 4455, 13 => 7151),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 19777, 3 => 6183, 4 => 9972, 5 => 14536, 6 => 8182, 7 => 17749, 8 => 11341, 9 => 5556, 10 => 4379, 11 => 17434, 12 => 15477, 13 => 18532),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 4651, 3 => 19689, 4 => 1608, 5 => 659, 6 => 16707, 7 => 14335, 8 => 6143, 9 => 3058, 10 => 14618, 11 => 17894, 12 => 20684, 13 => 5306),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 9778, 3 => 2552, 4 => 12096, 5 => 12369, 6 => 15198, 7 => 16890, 8 => 4851, 9 => 3109, 10 => 1700, 11 => 18725, 12 => 1997, 13 => 15882),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 486, 3 => 6111, 4 => 13743, 5 => 11537, 6 => 5591, 7 => 7433, 8 => 15227, 9 => 14145, 10 => 1483, 11 => 3887, 12 => 17431, 13 => 12430),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 20647, 3 => 14311, 4 => 11734, 5 => 4180, 6 => 8110, 7 => 5525, 8 => 12141, 9 => 15761, 10 => 18661, 11 => 18441, 12 => 10569, 13 => 8192),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 3791, 3 => 14759, 4 => 15264, 5 => 19918, 6 => 10132, 7 => 9062, 8 => 10010, 9 => 12786, 10 => 10675, 11 => 9682, 12 => 19246, 13 => 5454),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 19525, 3 => 9485, 4 => 7777, 5 => 19999, 6 => 8378, 7 => 9209, 8 => 3163, 9 => 20232, 10 => 6690, 11 => 16518, 12 => 716, 13 => 7353),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 4588, 3 => 6709, 4 => 20202, 5 => 10905, 6 => 915, 7 => 4317, 8 => 11073, 9 => 13576, 10 => 16433, 11 => 368, 12 => 3508, 13 => 21171),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 14072, 3 => 4033, 4 => 19959, 5 => 12608, 6 => 631, 7 => 19494, 8 => 14160, 9 => 8249, 10 => 10223, 11 => 21504, 12 => 12395, 13 => 4322),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 13800, 3 => 14161, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2948, 3 => 9647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 14693, 3 => 16027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 20506, 3 => 11082, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1143, 3 => 9020, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13501, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1548, 3 => 2190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 12216, 3 => 21556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 19897, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4189, 3 => 7958, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 15940, 3 => 10048, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 515, 3 => 12614, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8501, 3 => 8450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 17595, 3 => 16784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 5913, 3 => 8495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 16394, 3 => 10423, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7409, 3 => 6981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6678, 3 => 15939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20344, 3 => 12987, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 2510, 3 => 14588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 17918, 3 => 6655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 6703, 3 => 19451, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 496, 3 => 4217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7290, 3 => 5766, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 10521, 3 => 8925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 20379, 3 => 11905, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4090, 3 => 5838, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 19082, 3 => 17040, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 20233, 3 => 12352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 19365, 3 => 19546, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6249, 3 => 19030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11037, 3 => 19193, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 19760, 3 => 11772, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 45, 2 => 19644, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16076, 3 => 3521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11779, 3 => 21062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 48, 2 => 13062, 3 => 9682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 49, 2 => 8934, 3 => 5217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 50, 2 => 11087, 3 => 3319, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 51, 2 => 18892, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 52, 2 => 7894, 3 => 3898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 53, 2 => 5963, 3 => 4360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 54, 2 => 7346, 3 => 11726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5182, 3 => 5609, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 56, 2 => 2412, 3 => 17295, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 57, 2 => 9845, 3 => 20494, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 58, 2 => 6687, 3 => 1864, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 59, 2 => 20564, 3 => 5216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18226, 3 => 17207, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9380, 3 => 8266, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7073, 3 => 3065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 18252, 3 => 13437, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9161, 3 => 15642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10714, 3 => 10153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 11585, 3 => 9078, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5359, 3 => 9418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 9024, 3 => 9515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1206, 3 => 16354, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 14994, 3 => 1102, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9375, 3 => 20796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 15964, 3 => 6027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14789, 3 => 6452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8002, 3 => 18591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 14742, 3 => 14089, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 253, 3 => 3045, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1274, 3 => 19286, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 14777, 3 => 2044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 13920, 3 => 9900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 452, 3 => 7374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 18206, 3 => 9921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6131, 3 => 5414, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10077, 3 => 9726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 12045, 3 => 5479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4322, 3 => 7990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 15616, 3 => 5550, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 15561, 3 => 10661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 20718, 3 => 7387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2518, 3 => 18804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8984, 3 => 2600, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6516, 3 => 17909, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 32, 2 => 11148, 3 => 98, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 33, 2 => 20559, 3 => 3704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7510, 3 => 1569, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 35, 2 => 16000, 3 => 11692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 36, 2 => 9147, 3 => 10303, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 37, 2 => 16650, 3 => 191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15577, 3 => 18685, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 39, 2 => 17167, 3 => 20917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 40, 2 => 4256, 3 => 3391, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 41, 2 => 20092, 3 => 17219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 42, 2 => 9218, 3 => 5056, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 43, 2 => 18429, 3 => 8472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12093, 3 => 20753, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 45, 2 => 16345, 3 => 12748, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16023, 3 => 11095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 47, 2 => 5048, 3 => 17595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 48, 2 => 18995, 3 => 4817, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 49, 2 => 16483, 3 => 3536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 50, 2 => 1439, 3 => 16148, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 51, 2 => 3661, 3 => 3039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 52, 2 => 19010, 3 => 18121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 53, 2 => 8968, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 54, 2 => 13427, 3 => 18003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5303, 3 => 3083, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 56, 2 => 531, 3 => 16668, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 57, 2 => 4771, 3 => 6722, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 58, 2 => 5695, 3 => 7960, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 59, 2 => 3589, 3 => 14630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_5.csv, table is 72x196 (1764.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5 : integer_2d_array_t(0 to 71)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 31413, 2 => 18834, 3 => 28884, 4 => 947, 5 => 23050, 6 => 14484, 7 => 14809, 8 => 4968, 9 => 455, 10 => 33659, 11 => 16666, 12 => 19008),
    1 => integer_vector_t'(0 => 12, 1 => 13172, 2 => 19939, 3 => 13354, 4 => 13719, 5 => 6132, 6 => 20086, 7 => 34040, 8 => 13442, 9 => 27958, 10 => 16813, 11 => 29619, 12 => 16553),
    2 => integer_vector_t'(0 => 12, 1 => 1499, 2 => 32075, 3 => 14962, 4 => 11578, 5 => 11204, 6 => 9217, 7 => 10485, 8 => 23062, 9 => 30936, 10 => 17892, 11 => 24204, 12 => 24885),
    3 => integer_vector_t'(0 => 12, 1 => 32490, 2 => 18086, 3 => 18007, 4 => 4957, 5 => 7285, 6 => 32073, 7 => 19038, 8 => 7152, 9 => 12486, 10 => 13483, 11 => 24808, 12 => 21759),
    4 => integer_vector_t'(0 => 12, 1 => 32321, 2 => 10839, 3 => 15620, 4 => 33521, 5 => 23030, 6 => 10646, 7 => 26236, 8 => 19744, 9 => 21713, 10 => 36784, 11 => 8016, 12 => 12869),
    5 => integer_vector_t'(0 => 12, 1 => 35597, 2 => 11129, 3 => 17948, 4 => 26160, 5 => 14729, 6 => 31943, 7 => 20416, 8 => 10000, 9 => 7882, 10 => 31380, 11 => 27858, 12 => 33356),
    6 => integer_vector_t'(0 => 12, 1 => 14125, 2 => 12131, 3 => 36199, 4 => 4058, 5 => 35992, 6 => 36594, 7 => 33698, 8 => 15475, 9 => 1566, 10 => 18498, 11 => 12725, 12 => 7067),
    7 => integer_vector_t'(0 => 12, 1 => 17406, 2 => 8372, 3 => 35437, 4 => 2888, 5 => 1184, 6 => 30068, 7 => 25802, 8 => 11056, 9 => 5507, 10 => 26313, 11 => 32205, 12 => 37232),
    8 => integer_vector_t'(0 => 12, 1 => 15254, 2 => 5365, 3 => 17308, 4 => 22519, 5 => 35009, 6 => 718, 7 => 5240, 8 => 16778, 9 => 23131, 10 => 24092, 11 => 20587, 12 => 33385),
    9 => integer_vector_t'(0 => 12, 1 => 27455, 2 => 17602, 3 => 4590, 4 => 21767, 5 => 22266, 6 => 27357, 7 => 30400, 8 => 8732, 9 => 5596, 10 => 3060, 11 => 33703, 12 => 3596),
    10 => integer_vector_t'(0 => 12, 1 => 6882, 2 => 873, 3 => 10997, 4 => 24738, 5 => 20770, 6 => 10067, 7 => 13379, 8 => 27409, 9 => 25463, 10 => 2673, 11 => 6998, 12 => 31378),
    11 => integer_vector_t'(0 => 12, 1 => 15181, 2 => 13645, 3 => 34501, 4 => 3393, 5 => 3840, 6 => 35227, 7 => 15562, 8 => 23615, 9 => 38342, 10 => 12139, 11 => 19471, 12 => 15483),
    12 => integer_vector_t'(0 => 12, 1 => 13350, 2 => 6707, 3 => 23709, 4 => 37204, 5 => 25778, 6 => 21082, 7 => 7511, 8 => 14588, 9 => 10010, 10 => 21854, 11 => 28375, 12 => 33591),
    13 => integer_vector_t'(0 => 12, 1 => 12514, 2 => 4695, 3 => 37190, 4 => 21379, 5 => 18723, 6 => 5802, 7 => 7182, 8 => 2529, 9 => 29936, 10 => 35860, 11 => 28338, 12 => 10835),
    14 => integer_vector_t'(0 => 12, 1 => 34283, 2 => 25610, 3 => 33026, 4 => 31017, 5 => 21259, 6 => 2165, 7 => 21807, 8 => 37578, 9 => 1175, 10 => 16710, 11 => 21939, 12 => 30841),
    15 => integer_vector_t'(0 => 12, 1 => 27292, 2 => 33730, 3 => 6836, 4 => 26476, 5 => 27539, 6 => 35784, 7 => 18245, 8 => 16394, 9 => 17939, 10 => 23094, 11 => 19216, 12 => 17432),
    16 => integer_vector_t'(0 => 12, 1 => 11655, 2 => 6183, 3 => 38708, 4 => 28408, 5 => 35157, 6 => 17089, 7 => 13998, 8 => 36029, 9 => 15052, 10 => 16617, 11 => 5638, 12 => 36464),
    17 => integer_vector_t'(0 => 12, 1 => 15693, 2 => 28923, 3 => 26245, 4 => 9432, 5 => 11675, 6 => 25720, 7 => 26405, 8 => 5838, 9 => 31851, 10 => 26898, 11 => 8090, 12 => 37037),
    18 => integer_vector_t'(0 => 12, 1 => 24418, 2 => 27583, 3 => 7959, 4 => 35562, 5 => 37771, 6 => 17784, 7 => 11382, 8 => 11156, 9 => 37855, 10 => 7073, 11 => 21685, 12 => 34515),
    19 => integer_vector_t'(0 => 12, 1 => 10977, 2 => 13633, 3 => 30969, 4 => 7516, 5 => 11943, 6 => 18199, 7 => 5231, 8 => 13825, 9 => 19589, 10 => 23661, 11 => 11150, 12 => 35602),
    20 => integer_vector_t'(0 => 12, 1 => 19124, 2 => 30774, 3 => 6670, 4 => 37344, 5 => 16510, 6 => 26317, 7 => 23518, 8 => 22957, 9 => 6348, 10 => 34069, 11 => 8845, 12 => 20175),
    21 => integer_vector_t'(0 => 12, 1 => 34985, 2 => 14441, 3 => 25668, 4 => 4116, 5 => 3019, 6 => 21049, 7 => 37308, 8 => 24551, 9 => 24727, 10 => 20104, 11 => 24850, 12 => 12114),
    22 => integer_vector_t'(0 => 12, 1 => 38187, 2 => 28527, 3 => 13108, 4 => 13985, 5 => 1425, 6 => 21477, 7 => 30807, 8 => 8613, 9 => 26241, 10 => 33368, 11 => 35913, 12 => 32477),
    23 => integer_vector_t'(0 => 12, 1 => 5903, 2 => 34390, 3 => 24641, 4 => 26556, 5 => 23007, 6 => 27305, 7 => 38247, 8 => 2621, 9 => 9122, 10 => 32806, 11 => 21554, 12 => 18685),
    24 => integer_vector_t'(0 => 3, 1 => 17287, 2 => 27292, 3 => 19033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25796, 2 => 31795, 3 => 12152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 12184, 2 => 35088, 3 => 31226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 38263, 2 => 33386, 3 => 24892, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 23114, 2 => 37995, 3 => 29796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 34336, 2 => 10551, 3 => 36245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 35407, 2 => 175, 3 => 7203, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14654, 2 => 38201, 3 => 22605, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 28404, 2 => 6595, 3 => 1018, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 19932, 2 => 3524, 3 => 29305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 31749, 2 => 20247, 3 => 8128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 18026, 2 => 36357, 3 => 26735, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7543, 2 => 29767, 3 => 13588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 13333, 2 => 25965, 3 => 8463, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 14504, 2 => 36796, 3 => 19710, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4528, 2 => 25299, 3 => 7318, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 35091, 2 => 25550, 3 => 14798, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 7824, 2 => 215, 3 => 1248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 30848, 2 => 5362, 3 => 17291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 28932, 2 => 30249, 3 => 27073, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 13062, 2 => 2103, 3 => 16206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 7129, 2 => 32062, 3 => 19612, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 9512, 2 => 21936, 3 => 38833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 35849, 2 => 33754, 3 => 23450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18705, 2 => 28656, 3 => 18111, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 22749, 2 => 27456, 3 => 32187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 28229, 2 => 31684, 3 => 30160, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15293, 2 => 8483, 3 => 28002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 14880, 2 => 13334, 3 => 12584, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 28646, 2 => 2558, 3 => 19687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 6259, 2 => 4499, 3 => 26336, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 11952, 2 => 28386, 3 => 8405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 10609, 2 => 961, 3 => 7582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 10423, 2 => 13191, 3 => 26818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 15922, 2 => 36654, 3 => 21450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 10492, 2 => 1532, 3 => 1205, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 30551, 2 => 36482, 3 => 22153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 5156, 2 => 11330, 3 => 34243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 28616, 2 => 35369, 3 => 13322, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 8962, 2 => 1485, 3 => 21186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 23541, 2 => 17445, 3 => 35561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 33133, 2 => 11593, 3 => 19895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 33917, 2 => 7863, 3 => 33651, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 20063, 2 => 28331, 3 => 10702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 13195, 2 => 21107, 3 => 21859, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 4364, 2 => 31137, 3 => 4804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 5585, 2 => 2037, 3 => 4830, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 30672, 2 => 16927, 3 => 14800, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_4.csv, table is 135x164 (2767.5 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4 : integer_2d_array_t(0 to 134)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 0, 2 => 6385, 3 => 7901, 4 => 14611, 5 => 13389, 6 => 11200, 7 => 3252, 8 => 5243, 9 => 2504, 10 => 2722, 11 => 821, 12 => 7374),
    1 => integer_vector_t'(0 => 12, 1 => 1, 2 => 11359, 3 => 2698, 4 => 357, 5 => 13824, 6 => 12772, 7 => 7244, 8 => 6752, 9 => 15310, 10 => 852, 11 => 2001, 12 => 11417),
    2 => integer_vector_t'(0 => 12, 1 => 2, 2 => 7862, 3 => 7977, 4 => 6321, 5 => 13612, 6 => 12197, 7 => 14449, 8 => 15137, 9 => 13860, 10 => 1708, 11 => 6399, 12 => 13444),
    3 => integer_vector_t'(0 => 12, 1 => 3, 2 => 1560, 3 => 11804, 4 => 6975, 5 => 13292, 6 => 3646, 7 => 3812, 8 => 8772, 9 => 7306, 10 => 5795, 11 => 14327, 12 => 7866),
    4 => integer_vector_t'(0 => 12, 1 => 4, 2 => 7626, 3 => 11407, 4 => 14599, 5 => 9689, 6 => 1628, 7 => 2113, 8 => 10809, 9 => 9283, 10 => 1230, 11 => 15241, 12 => 4870),
    5 => integer_vector_t'(0 => 12, 1 => 5, 2 => 1610, 3 => 5699, 4 => 15876, 5 => 9446, 6 => 12515, 7 => 1400, 8 => 6303, 9 => 5411, 10 => 14181, 11 => 13925, 12 => 7358),
    6 => integer_vector_t'(0 => 12, 1 => 6, 2 => 4059, 3 => 8836, 4 => 3405, 5 => 7853, 6 => 7992, 7 => 15336, 8 => 5970, 9 => 10368, 10 => 10278, 11 => 9675, 12 => 4651),
    7 => integer_vector_t'(0 => 12, 1 => 7, 2 => 4441, 3 => 3963, 4 => 9153, 5 => 2109, 6 => 12683, 7 => 7459, 8 => 12030, 9 => 12221, 10 => 629, 11 => 15212, 12 => 406),
    8 => integer_vector_t'(0 => 12, 1 => 8, 2 => 6007, 3 => 8411, 4 => 5771, 5 => 3497, 6 => 543, 7 => 14202, 8 => 875, 9 => 9186, 10 => 6235, 11 => 13908, 12 => 3563),
    9 => integer_vector_t'(0 => 12, 1 => 9, 2 => 3232, 3 => 6625, 4 => 4795, 5 => 546, 6 => 9781, 7 => 2071, 8 => 7312, 9 => 3399, 10 => 7250, 11 => 4932, 12 => 12652),
    10 => integer_vector_t'(0 => 12, 1 => 10, 2 => 8820, 3 => 10088, 4 => 11090, 5 => 7069, 6 => 6585, 7 => 13134, 8 => 10158, 9 => 7183, 10 => 488, 11 => 7455, 12 => 9238),
    11 => integer_vector_t'(0 => 12, 1 => 11, 2 => 1903, 3 => 10818, 4 => 119, 5 => 215, 6 => 7558, 7 => 11046, 8 => 10615, 9 => 11545, 10 => 14784, 11 => 7961, 12 => 15619),
    12 => integer_vector_t'(0 => 12, 1 => 12, 2 => 3655, 3 => 8736, 4 => 4917, 5 => 15874, 6 => 5129, 7 => 2134, 8 => 15944, 9 => 14768, 10 => 7150, 11 => 2692, 12 => 1469),
    13 => integer_vector_t'(0 => 12, 1 => 13, 2 => 8316, 3 => 3820, 4 => 505, 5 => 8923, 6 => 6757, 7 => 806, 8 => 7957, 9 => 4216, 10 => 15589, 11 => 13244, 12 => 2622),
    14 => integer_vector_t'(0 => 12, 1 => 14, 2 => 14463, 3 => 4852, 4 => 15733, 5 => 3041, 6 => 11193, 7 => 12860, 8 => 13673, 9 => 8152, 10 => 6551, 11 => 15108, 12 => 8758),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3149, 3 => 11981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 13416, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13098, 3 => 13352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 2009, 3 => 14460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 7207, 3 => 4314, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 3312, 3 => 3945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4418, 3 => 6248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 2669, 3 => 13975, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 7571, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14172, 3 => 2967, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7271, 3 => 7138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6135, 3 => 13670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 7490, 3 => 14559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8657, 3 => 2466, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8599, 3 => 12834, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 3470, 3 => 3152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13917, 3 => 4365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 6024, 3 => 13730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 10973, 3 => 14182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 2464, 3 => 13167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 5281, 3 => 15049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 1103, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 2058, 3 => 1069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 9654, 3 => 6095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 14311, 3 => 7667, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 15617, 3 => 8146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 4588, 3 => 11218, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 13660, 3 => 6243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 8578, 3 => 7874, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 11741, 3 => 2686, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1022, 3 => 1264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 1, 2 => 12604, 3 => 9965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 2, 2 => 8217, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3156, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 4, 2 => 354, 3 => 1514, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6978, 3 => 14058, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 6, 2 => 7922, 3 => 16079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 7, 2 => 15087, 3 => 12138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5053, 3 => 6470, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 9, 2 => 12687, 3 => 14932, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15458, 3 => 1763, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8121, 3 => 1721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 12, 2 => 12431, 3 => 549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4129, 3 => 7091, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1426, 3 => 8415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9783, 3 => 7604, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6295, 3 => 11329, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1409, 3 => 12061, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 18, 2 => 8065, 3 => 9087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2918, 3 => 8438, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1293, 3 => 14115, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 21, 2 => 3922, 3 => 13851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3851, 3 => 4000, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5865, 3 => 1768, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2655, 3 => 14957, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 25, 2 => 5565, 3 => 6332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4303, 3 => 12631, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11653, 3 => 12236, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 28, 2 => 16025, 3 => 7632, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4655, 3 => 14128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 30, 2 => 9584, 3 => 13123, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13987, 3 => 9597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 32, 2 => 15409, 3 => 12110, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 33, 2 => 8754, 3 => 15490, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7416, 3 => 15325, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2909, 3 => 15549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 36, 2 => 2995, 3 => 8257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 37, 2 => 9406, 3 => 4791, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 38, 2 => 11111, 3 => 4854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 39, 2 => 2812, 3 => 8521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 40, 2 => 8476, 3 => 14717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7820, 3 => 15360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 42, 2 => 1179, 3 => 7939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 43, 2 => 2357, 3 => 8678, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 44, 2 => 7703, 3 => 6216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3477, 3 => 7067, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3931, 3 => 13845, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7675, 3 => 12899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1754, 3 => 8187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7785, 3 => 1400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 9213, 3 => 5891, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2494, 3 => 7703, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2576, 3 => 7902, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4821, 3 => 15682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 10426, 3 => 11935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1810, 3 => 904, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 11332, 3 => 9264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11312, 3 => 3570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14916, 3 => 2650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7679, 3 => 7842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6089, 3 => 13084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3938, 3 => 2751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8509, 3 => 4648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 12204, 3 => 8917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5749, 3 => 12443, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12613, 3 => 4431, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1344, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 8488, 3 => 13850, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1730, 3 => 14896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14942, 3 => 7126, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 14983, 3 => 8863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6578, 3 => 8564, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 4947, 3 => 396, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 297, 3 => 12805, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 13878, 3 => 6692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11857, 3 => 11186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 31, 2 => 14395, 3 => 11493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 32, 2 => 16145, 3 => 12251, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 33, 2 => 13462, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 34, 2 => 14526, 3 => 13119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2535, 3 => 11243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 36, 2 => 6465, 3 => 12690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 37, 2 => 6872, 3 => 9334, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15371, 3 => 14023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 39, 2 => 8101, 3 => 10187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 40, 2 => 11963, 3 => 4848, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 41, 2 => 15125, 3 => 6119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 42, 2 => 8051, 3 => 14465, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11139, 3 => 5167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 44, 2 => 2883, 3 => 14521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_5.csv, table is 108x184 (2484.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 15, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15, 9 => 15, 10 => 15, 11 => 15, 12 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5 : integer_2d_array_t(0 to 107)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 22422, 2 => 10282, 3 => 11626, 4 => 19997, 5 => 11161, 6 => 2922, 7 => 3122, 8 => 99, 9 => 5625, 10 => 17064, 11 => 8270, 12 => 179),
    1 => integer_vector_t'(0 => 12, 1 => 25087, 2 => 16218, 3 => 17015, 4 => 828, 5 => 20041, 6 => 25656, 7 => 4186, 8 => 11629, 9 => 22599, 10 => 17305, 11 => 22515, 12 => 6463),
    2 => integer_vector_t'(0 => 12, 1 => 11049, 2 => 22853, 3 => 25706, 4 => 14388, 5 => 5500, 6 => 19245, 7 => 8732, 8 => 2177, 9 => 13555, 10 => 11346, 11 => 17265, 12 => 3069),
    3 => integer_vector_t'(0 => 12, 1 => 16581, 2 => 22225, 3 => 12563, 4 => 19717, 5 => 23577, 6 => 11555, 7 => 25496, 8 => 6853, 9 => 25403, 10 => 5218, 11 => 15925, 12 => 21766),
    4 => integer_vector_t'(0 => 12, 1 => 16529, 2 => 14487, 3 => 7643, 4 => 10715, 5 => 17442, 6 => 11119, 7 => 5679, 8 => 14155, 9 => 24213, 10 => 21000, 11 => 1116, 12 => 15620),
    5 => integer_vector_t'(0 => 12, 1 => 5340, 2 => 8636, 3 => 16693, 4 => 1434, 5 => 5635, 6 => 6516, 7 => 9482, 8 => 20189, 9 => 1066, 10 => 15013, 11 => 25361, 12 => 14243),
    6 => integer_vector_t'(0 => 12, 1 => 18506, 2 => 22236, 3 => 20912, 4 => 8952, 5 => 5421, 6 => 15691, 7 => 6126, 8 => 21595, 9 => 500, 10 => 6904, 11 => 13059, 12 => 6802),
    7 => integer_vector_t'(0 => 12, 1 => 8433, 2 => 4694, 3 => 5524, 4 => 14216, 5 => 3685, 6 => 19721, 7 => 25420, 8 => 9937, 9 => 23813, 10 => 9047, 11 => 25651, 12 => 16826),
    8 => integer_vector_t'(0 => 12, 1 => 21500, 2 => 24814, 3 => 6344, 4 => 17382, 5 => 7064, 6 => 13929, 7 => 4004, 8 => 16552, 9 => 12818, 10 => 8720, 11 => 5286, 12 => 2206),
    9 => integer_vector_t'(0 => 12, 1 => 22517, 2 => 2429, 3 => 19065, 4 => 2921, 5 => 21611, 6 => 1873, 7 => 7507, 8 => 5661, 9 => 23006, 10 => 23128, 11 => 20543, 12 => 19777),
    10 => integer_vector_t'(0 => 12, 1 => 1770, 2 => 4636, 3 => 20900, 4 => 14931, 5 => 9247, 6 => 12340, 7 => 11008, 8 => 12966, 9 => 4471, 10 => 2731, 11 => 16445, 12 => 791),
    11 => integer_vector_t'(0 => 12, 1 => 6635, 2 => 14556, 3 => 18865, 4 => 22421, 5 => 22124, 6 => 12697, 7 => 9803, 8 => 25485, 9 => 7744, 10 => 18254, 11 => 11313, 12 => 9004),
    12 => integer_vector_t'(0 => 12, 1 => 19982, 2 => 23963, 3 => 18912, 4 => 7206, 5 => 12500, 6 => 4382, 7 => 20067, 8 => 6177, 9 => 21007, 10 => 1195, 11 => 23547, 12 => 24837),
    13 => integer_vector_t'(0 => 12, 1 => 756, 2 => 11158, 3 => 14646, 4 => 20534, 5 => 3647, 6 => 17728, 7 => 11676, 8 => 11843, 9 => 12937, 10 => 4402, 11 => 8261, 12 => 22944),
    14 => integer_vector_t'(0 => 12, 1 => 9306, 2 => 24009, 3 => 10012, 4 => 11081, 5 => 3746, 6 => 24325, 7 => 8060, 8 => 19826, 9 => 842, 10 => 8836, 11 => 2898, 12 => 5019),
    15 => integer_vector_t'(0 => 12, 1 => 7575, 2 => 7455, 3 => 25244, 4 => 4736, 5 => 14400, 6 => 22981, 7 => 5543, 8 => 8006, 9 => 24203, 10 => 13053, 11 => 1120, 12 => 5128),
    16 => integer_vector_t'(0 => 12, 1 => 3482, 2 => 9270, 3 => 13059, 4 => 15825, 5 => 7453, 6 => 23747, 7 => 3656, 8 => 24585, 9 => 16542, 10 => 17507, 11 => 22462, 12 => 14670),
    17 => integer_vector_t'(0 => 12, 1 => 15627, 2 => 15290, 3 => 4198, 4 => 22748, 5 => 5842, 6 => 13395, 7 => 23918, 8 => 16985, 9 => 14929, 10 => 3726, 11 => 25350, 12 => 24157),
    18 => integer_vector_t'(0 => 12, 1 => 24896, 2 => 16365, 3 => 16423, 4 => 13461, 5 => 16615, 6 => 8107, 7 => 24741, 8 => 3604, 9 => 25904, 10 => 8716, 11 => 9604, 12 => 20365),
    19 => integer_vector_t'(0 => 12, 1 => 3729, 2 => 17245, 3 => 18448, 4 => 9862, 5 => 20831, 6 => 25326, 7 => 20517, 8 => 24618, 9 => 13282, 10 => 5099, 11 => 14183, 12 => 8804),
    20 => integer_vector_t'(0 => 12, 1 => 16455, 2 => 17646, 3 => 15376, 4 => 18194, 5 => 25528, 6 => 1777, 7 => 6066, 8 => 21855, 9 => 14372, 10 => 12517, 11 => 4488, 12 => 17490),
    21 => integer_vector_t'(0 => 12, 1 => 1400, 2 => 8135, 3 => 23375, 4 => 20879, 5 => 8476, 6 => 4084, 7 => 12936, 8 => 25536, 9 => 22309, 10 => 16582, 11 => 6402, 12 => 24360),
    22 => integer_vector_t'(0 => 12, 1 => 25119, 2 => 23586, 3 => 128, 4 => 4761, 5 => 10443, 6 => 22536, 7 => 8607, 8 => 9752, 9 => 25446, 10 => 15053, 11 => 1856, 12 => 4040),
    23 => integer_vector_t'(0 => 12, 1 => 377, 2 => 21160, 3 => 13474, 4 => 5451, 5 => 17170, 6 => 5938, 7 => 10256, 8 => 11972, 9 => 24210, 10 => 17833, 11 => 22047, 12 => 16108),
    24 => integer_vector_t'(0 => 12, 1 => 13075, 2 => 9648, 3 => 24546, 4 => 13150, 5 => 23867, 6 => 7309, 7 => 19798, 8 => 2988, 9 => 16858, 10 => 4825, 11 => 23950, 12 => 15125),
    25 => integer_vector_t'(0 => 12, 1 => 20526, 2 => 3553, 3 => 11525, 4 => 23366, 5 => 2452, 6 => 17626, 7 => 19265, 8 => 20172, 9 => 18060, 10 => 24593, 11 => 13255, 12 => 1552),
    26 => integer_vector_t'(0 => 12, 1 => 18839, 2 => 21132, 3 => 20119, 4 => 15214, 5 => 14705, 6 => 7096, 7 => 10174, 8 => 5663, 9 => 18651, 10 => 19700, 11 => 12524, 12 => 14033),
    27 => integer_vector_t'(0 => 12, 1 => 4127, 2 => 2971, 3 => 17499, 4 => 16287, 5 => 22368, 6 => 21463, 7 => 7943, 8 => 18880, 9 => 5567, 10 => 8047, 11 => 23363, 12 => 6797),
    28 => integer_vector_t'(0 => 12, 1 => 10651, 2 => 24471, 3 => 14325, 4 => 4081, 5 => 7258, 6 => 4949, 7 => 7044, 8 => 1078, 9 => 797, 10 => 22910, 11 => 20474, 12 => 4318),
    29 => integer_vector_t'(0 => 12, 1 => 21374, 2 => 13231, 3 => 22985, 4 => 5056, 5 => 3821, 6 => 23718, 7 => 14178, 8 => 9978, 9 => 19030, 10 => 23594, 11 => 8895, 12 => 25358),
    30 => integer_vector_t'(0 => 12, 1 => 6199, 2 => 22056, 3 => 7749, 4 => 13310, 5 => 3999, 6 => 23697, 7 => 16445, 8 => 22636, 9 => 5225, 10 => 22437, 11 => 24153, 12 => 9442),
    31 => integer_vector_t'(0 => 12, 1 => 7978, 2 => 12177, 3 => 2893, 4 => 20778, 5 => 3175, 6 => 8645, 7 => 11863, 8 => 24623, 9 => 10311, 10 => 25767, 11 => 17057, 12 => 3691),
    32 => integer_vector_t'(0 => 12, 1 => 20473, 2 => 11294, 3 => 9914, 4 => 22815, 5 => 2574, 6 => 8439, 7 => 3699, 8 => 5431, 9 => 24840, 10 => 21908, 11 => 16088, 12 => 18244),
    33 => integer_vector_t'(0 => 12, 1 => 8208, 2 => 5755, 3 => 19059, 4 => 8541, 5 => 24924, 6 => 6454, 7 => 11234, 8 => 10492, 9 => 16406, 10 => 10831, 11 => 11436, 12 => 9649),
    34 => integer_vector_t'(0 => 12, 1 => 16264, 2 => 11275, 3 => 24953, 4 => 2347, 5 => 12667, 6 => 19190, 7 => 7257, 8 => 7174, 9 => 24819, 10 => 2938, 11 => 2522, 12 => 11749),
    35 => integer_vector_t'(0 => 12, 1 => 3627, 2 => 5969, 3 => 13862, 4 => 1538, 5 => 23176, 6 => 6353, 7 => 2855, 8 => 17720, 9 => 2472, 10 => 7428, 11 => 573, 12 => 15036),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18539, 3 => 18661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 10502, 3 => 3002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 9368, 3 => 10761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 12299, 3 => 7828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 15048, 3 => 13362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 18444, 3 => 24640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 20775, 3 => 19175, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 18970, 3 => 10971, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5329, 3 => 19982, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 11296, 3 => 18655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15046, 3 => 20659, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 7300, 3 => 22140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 22029, 3 => 14477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 11129, 3 => 742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 13254, 3 => 13813, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 19234, 3 => 13273, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6079, 3 => 21122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 22782, 3 => 5828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 19775, 3 => 4247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1660, 3 => 19413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4403, 3 => 3649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 13371, 3 => 25851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 22770, 3 => 21784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10757, 3 => 14131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 16071, 3 => 21617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 6393, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 597, 3 => 19968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5743, 3 => 8084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 6770, 3 => 9548, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4285, 3 => 17542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 13568, 3 => 22599, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 1786, 3 => 4617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 23238, 3 => 11648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 19627, 3 => 2030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 13601, 3 => 13458, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 13740, 3 => 17328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 25012, 3 => 13944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 22513, 3 => 6687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4934, 3 => 12587, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 21197, 3 => 5133, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 22705, 3 => 6938, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7534, 3 => 24633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 24400, 3 => 12797, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 21911, 3 => 25712, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12039, 3 => 1140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 24306, 3 => 1021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 14012, 3 => 20747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11265, 3 => 15219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 4670, 3 => 15531, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 9417, 3 => 14359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 2415, 3 => 6504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 24964, 3 => 24690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 14443, 3 => 8816, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 6926, 3 => 1291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 54, 2 => 6209, 3 => 20806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 55, 2 => 13915, 3 => 4079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 56, 2 => 24410, 3 => 13196, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 57, 2 => 13505, 3 => 6117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 58, 2 => 9869, 3 => 8220, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 59, 2 => 1570, 3 => 6044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 60, 2 => 25780, 3 => 17387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 61, 2 => 20671, 3 => 24913, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 62, 2 => 24558, 3 => 20591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 63, 2 => 12402, 3 => 3702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 64, 2 => 8314, 3 => 1357, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 65, 2 => 20071, 3 => 14616, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 66, 2 => 17014, 3 => 3688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 67, 2 => 19837, 3 => 946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 68, 2 => 15195, 3 => 12136, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 69, 2 => 7758, 3 => 22808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 70, 2 => 3564, 3 => 2925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 71, 2 => 3434, 3 => 7769, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C4_5.csv, table is 144x150 (2700.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5 : integer_2d_array_t(0 to 143)(0 to 11) := (
    0 => integer_vector_t'(0 => 11, 1 => 0, 2 => 149, 3 => 11212, 4 => 5575, 5 => 6360, 6 => 12559, 7 => 8108, 8 => 8505, 9 => 408, 10 => 10026, 11 => 12828),
    1 => integer_vector_t'(0 => 11, 1 => 1, 2 => 5237, 3 => 490, 4 => 10677, 5 => 4998, 6 => 3869, 7 => 3734, 8 => 3092, 9 => 3509, 10 => 7703, 11 => 10305),
    2 => integer_vector_t'(0 => 11, 1 => 2, 2 => 8742, 3 => 5553, 4 => 2820, 5 => 7085, 6 => 12116, 7 => 10485, 8 => 564, 9 => 7795, 10 => 2972, 11 => 2157),
    3 => integer_vector_t'(0 => 11, 1 => 3, 2 => 2699, 3 => 4304, 4 => 8350, 5 => 712, 6 => 2841, 7 => 3250, 8 => 4731, 9 => 10105, 10 => 517, 11 => 7516),
    4 => integer_vector_t'(0 => 11, 1 => 4, 2 => 12067, 3 => 1351, 4 => 11992, 5 => 12191, 6 => 11267, 7 => 5161, 8 => 537, 9 => 6166, 10 => 4246, 11 => 2363),
    5 => integer_vector_t'(0 => 11, 1 => 5, 2 => 6828, 3 => 7107, 4 => 2127, 5 => 3724, 6 => 5743, 7 => 11040, 8 => 10756, 9 => 4073, 10 => 1011, 11 => 3422),
    6 => integer_vector_t'(0 => 11, 1 => 6, 2 => 11259, 3 => 1216, 4 => 9526, 5 => 1466, 6 => 10816, 7 => 940, 8 => 3744, 9 => 2815, 10 => 11506, 11 => 11573),
    7 => integer_vector_t'(0 => 11, 1 => 7, 2 => 4549, 3 => 11507, 4 => 1118, 5 => 1274, 6 => 11751, 7 => 5207, 8 => 7854, 9 => 12803, 10 => 4047, 11 => 6484),
    8 => integer_vector_t'(0 => 11, 1 => 8, 2 => 8430, 3 => 4115, 4 => 9440, 5 => 413, 6 => 4455, 7 => 2262, 8 => 7915, 9 => 12402, 10 => 8579, 11 => 7052),
    9 => integer_vector_t'(0 => 11, 1 => 9, 2 => 3885, 3 => 9126, 4 => 5665, 5 => 4505, 6 => 2343, 7 => 253, 8 => 4707, 9 => 3742, 10 => 4166, 11 => 1556),
    10 => integer_vector_t'(0 => 11, 1 => 10, 2 => 1704, 3 => 8936, 4 => 6775, 5 => 8639, 6 => 8179, 7 => 7954, 8 => 8234, 9 => 7850, 10 => 8883, 11 => 8713),
    11 => integer_vector_t'(0 => 11, 1 => 11, 2 => 11716, 3 => 4344, 4 => 9087, 5 => 11264, 6 => 2274, 7 => 8832, 8 => 9147, 9 => 11930, 10 => 6054, 11 => 5455),
    12 => integer_vector_t'(0 => 11, 1 => 12, 2 => 7323, 3 => 3970, 4 => 10329, 5 => 2170, 6 => 8262, 7 => 3854, 8 => 2087, 9 => 12899, 10 => 9497, 11 => 11700),
    13 => integer_vector_t'(0 => 11, 1 => 13, 2 => 4418, 3 => 1467, 4 => 2490, 5 => 5841, 6 => 817, 7 => 11453, 8 => 533, 9 => 11217, 10 => 11962, 11 => 5251),
    14 => integer_vector_t'(0 => 11, 1 => 14, 2 => 1541, 3 => 4525, 4 => 7976, 5 => 3457, 6 => 9536, 7 => 7725, 8 => 3788, 9 => 2982, 10 => 6307, 11 => 5997),
    15 => integer_vector_t'(0 => 11, 1 => 15, 2 => 11484, 3 => 2739, 4 => 4023, 5 => 12107, 6 => 6516, 7 => 551, 8 => 2572, 9 => 6628, 10 => 8150, 11 => 9852),
    16 => integer_vector_t'(0 => 11, 1 => 16, 2 => 6070, 3 => 1761, 4 => 4627, 5 => 6534, 6 => 7913, 7 => 3730, 8 => 11866, 9 => 1813, 10 => 12306, 11 => 8249),
    17 => integer_vector_t'(0 => 11, 1 => 17, 2 => 12441, 3 => 5489, 4 => 8748, 5 => 7837, 6 => 7660, 7 => 2102, 8 => 11341, 9 => 2936, 10 => 6712, 11 => 11977),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10155, 3 => 4210, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1010, 3 => 10483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 8900, 3 => 10250, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 10243, 3 => 12278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 7070, 3 => 4397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 12271, 3 => 3887, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 11980, 3 => 6836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 9514, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 7137, 3 => 10281, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11881, 3 => 2526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 1969, 3 => 11477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3044, 3 => 10921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 2236, 3 => 8724, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9104, 3 => 6340, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 7342, 3 => 8582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 11675, 3 => 10405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 6467, 3 => 12775, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 3186, 3 => 12198, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 9621, 3 => 11445, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7486, 3 => 5611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4319, 3 => 4879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2196, 3 => 344, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7527, 3 => 6650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10693, 3 => 2440, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6755, 3 => 2706, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5144, 3 => 5998, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 11043, 3 => 8033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4846, 3 => 4435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4157, 3 => 9228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 12270, 3 => 6562, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11954, 3 => 7592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 7420, 3 => 2592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8810, 3 => 9636, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 689, 3 => 5430, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 920, 3 => 1304, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1253, 3 => 11934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9559, 3 => 6016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 312, 3 => 7589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4439, 3 => 4197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4002, 3 => 9555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12232, 3 => 7779, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1494, 3 => 8782, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 10749, 3 => 3969, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4368, 3 => 3479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6316, 3 => 5342, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2455, 3 => 3493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12157, 3 => 7405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6598, 3 => 11495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11805, 3 => 4455, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9625, 3 => 2090, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 4731, 3 => 2321, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 3578, 3 => 2608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 8504, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 4027, 3 => 1151, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5647, 3 => 4935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4219, 3 => 1870, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10968, 3 => 8054, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6970, 3 => 5447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3217, 3 => 5638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 8972, 3 => 669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5618, 3 => 12472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1457, 3 => 1280, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 8868, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8866, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 8371, 3 => 5972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 266, 3 => 4405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3706, 3 => 3244, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 6039, 3 => 5844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7200, 3 => 3283, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1502, 3 => 11282, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 12318, 3 => 2202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4523, 3 => 965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9587, 3 => 7011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2552, 3 => 2051, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12045, 3 => 10306, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 21, 2 => 11070, 3 => 5104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6627, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 23, 2 => 9889, 3 => 2121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 24, 2 => 829, 3 => 9701, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2201, 3 => 1819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6689, 3 => 12925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2139, 3 => 8757, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12004, 3 => 5948, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8704, 3 => 3191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8171, 3 => 10933, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6297, 3 => 7116, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 32, 2 => 616, 3 => 7146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 33, 2 => 5142, 3 => 9761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 34, 2 => 10377, 3 => 8138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7616, 3 => 5811, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7285, 3 => 9863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7764, 3 => 10867, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 12343, 3 => 9019, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4414, 3 => 8331, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3464, 3 => 642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6960, 3 => 2039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 786, 3 => 3021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 710, 3 => 2086, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 7423, 3 => 5601, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8120, 3 => 4885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 12385, 3 => 11990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9739, 3 => 10034, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 424, 3 => 10162, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1347, 3 => 7597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1450, 3 => 112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 7965, 3 => 8478, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8945, 3 => 7397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 6590, 3 => 8316, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6838, 3 => 9011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6174, 3 => 9410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 20, 2 => 255, 3 => 113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 21, 2 => 6197, 3 => 5835, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12902, 3 => 3844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 23, 2 => 4377, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 24, 2 => 5478, 3 => 8672, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4453, 3 => 2132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 26, 2 => 9724, 3 => 1380, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 27, 2 => 12131, 3 => 11526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12323, 3 => 9511, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8231, 3 => 1752, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 30, 2 => 497, 3 => 9022, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9288, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 32, 2 => 2481, 3 => 7515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 33, 2 => 2696, 3 => 268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 34, 2 => 4023, 3 => 12341, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7108, 3 => 5553, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C5_6.csv, table is 150x177 (3318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 5, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14, 13 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6 : integer_2d_array_t(0 to 149)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 4362, 3 => 416, 4 => 8909, 5 => 4156, 6 => 3216, 7 => 3112, 8 => 2560, 9 => 2912, 10 => 6405, 11 => 8593, 12 => 4969, 13 => 6723),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 2479, 3 => 1786, 4 => 8978, 5 => 3011, 6 => 4339, 7 => 9313, 8 => 6397, 9 => 2957, 10 => 7288, 11 => 5484, 12 => 6031, 13 => 10217),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 10175, 3 => 9009, 4 => 9889, 5 => 3091, 6 => 4985, 7 => 7267, 8 => 4092, 9 => 8874, 10 => 5671, 11 => 2777, 12 => 2189, 13 => 8716),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 9052, 3 => 4795, 4 => 3924, 5 => 3370, 6 => 10058, 7 => 1128, 8 => 9996, 9 => 10165, 10 => 9360, 11 => 4297, 12 => 434, 13 => 5138),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 2379, 3 => 7834, 4 => 4835, 5 => 2327, 6 => 9843, 7 => 804, 8 => 329, 9 => 8353, 10 => 7167, 11 => 3070, 12 => 1528, 13 => 7311),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 3435, 3 => 7871, 4 => 348, 5 => 3693, 6 => 1876, 7 => 6585, 8 => 10340, 9 => 7144, 10 => 5870, 11 => 2084, 12 => 4052, 13 => 2780),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 3917, 3 => 3111, 4 => 3476, 5 => 1304, 6 => 10331, 7 => 5939, 8 => 5199, 9 => 1611, 10 => 1991, 11 => 699, 12 => 8316, 13 => 9960),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 6883, 3 => 3237, 4 => 1717, 5 => 10752, 6 => 7891, 7 => 9764, 8 => 4745, 9 => 3888, 10 => 10009, 11 => 4176, 12 => 4614, 13 => 1567),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 10587, 3 => 2195, 4 => 1689, 5 => 2968, 6 => 5420, 7 => 2580, 8 => 2883, 9 => 6496, 10 => 111, 11 => 6023, 12 => 1024, 13 => 4449),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 3786, 3 => 8593, 4 => 2074, 5 => 3321, 6 => 5057, 7 => 1450, 8 => 3840, 9 => 5444, 10 => 6572, 11 => 3094, 12 => 9892, 13 => 1512),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 8548, 3 => 1848, 4 => 10372, 5 => 4585, 6 => 7313, 7 => 6536, 8 => 6379, 9 => 1766, 10 => 9462, 11 => 2456, 12 => 5606, 13 => 9975),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 8204, 3 => 10593, 4 => 7935, 5 => 3636, 6 => 3882, 7 => 394, 8 => 5968, 9 => 8561, 10 => 2395, 11 => 7289, 12 => 9267, 13 => 9978),
    12 => integer_vector_t'(0 => 13, 1 => 12, 2 => 7795, 3 => 74, 4 => 1633, 5 => 9542, 6 => 6867, 7 => 7352, 8 => 6417, 9 => 7568, 10 => 10623, 11 => 725, 12 => 2531, 13 => 9115),
    13 => integer_vector_t'(0 => 13, 1 => 13, 2 => 7151, 3 => 2482, 4 => 4260, 5 => 5003, 6 => 10105, 7 => 7419, 8 => 9203, 9 => 6691, 10 => 8798, 11 => 2092, 12 => 8263, 13 => 3755),
    14 => integer_vector_t'(0 => 13, 1 => 14, 2 => 3600, 3 => 570, 4 => 4527, 5 => 200, 6 => 9718, 7 => 6771, 8 => 1995, 9 => 8902, 10 => 5446, 11 => 768, 12 => 1103, 13 => 6520),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6304, 3 => 7621, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6498, 3 => 9209, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 7293, 3 => 6786, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5950, 3 => 1708, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8521, 3 => 1793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 6174, 3 => 7854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9773, 3 => 1190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9517, 3 => 10268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2181, 3 => 9349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 1949, 3 => 5560, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 1556, 3 => 555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8600, 3 => 3827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5072, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7928, 3 => 3542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3226, 3 => 3762, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7045, 3 => 2420, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9645, 3 => 2641, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2774, 3 => 2452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5331, 3 => 2031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9400, 3 => 7503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1850, 3 => 2338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10456, 3 => 9774, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1692, 3 => 9276, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 8, 2 => 10037, 3 => 4038, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3964, 3 => 338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 10, 2 => 2640, 3 => 5087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 11, 2 => 858, 3 => 3473, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5582, 3 => 5683, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9523, 3 => 916, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4107, 3 => 1559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4506, 3 => 3491, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8191, 3 => 4182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 17, 2 => 10192, 3 => 6157, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5668, 3 => 3305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3449, 3 => 1540, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4766, 3 => 2697, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4069, 3 => 6675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 22, 2 => 1117, 3 => 1016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5619, 3 => 3085, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8483, 3 => 8400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 25, 2 => 8255, 3 => 394, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6338, 3 => 5042, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 27, 2 => 6174, 3 => 5119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7203, 3 => 1989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 29, 2 => 1781, 3 => 5174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1464, 3 => 3559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3376, 3 => 4214, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7238, 3 => 67, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 10595, 3 => 8831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1221, 3 => 6513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5300, 3 => 4652, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1429, 3 => 9749, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7878, 3 => 5131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4435, 3 => 10284, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6331, 3 => 5507, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6662, 3 => 4941, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9614, 3 => 10238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 8400, 3 => 8025, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9156, 3 => 5630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7067, 3 => 8878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9027, 3 => 3415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1690, 3 => 3866, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2854, 3 => 8469, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6206, 3 => 630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 363, 3 => 5453, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4125, 3 => 7008, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1612, 3 => 6702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9069, 3 => 9226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5767, 3 => 4060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 3743, 3 => 9237, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7018, 3 => 5572, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8892, 3 => 4536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 853, 3 => 6064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8069, 3 => 5893, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2051, 3 => 2885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 10691, 3 => 3153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3602, 3 => 4055, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 328, 3 => 1717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2219, 3 => 9299, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1939, 3 => 7898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 617, 3 => 206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 8544, 3 => 1374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 10676, 3 => 3240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6672, 3 => 9489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3170, 3 => 7457, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7868, 3 => 5731, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6121, 3 => 10732, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4843, 3 => 9132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 580, 3 => 9591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 6267, 3 => 9290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3009, 3 => 2268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 195, 3 => 2419, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8016, 3 => 1557, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1516, 3 => 9195, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8062, 3 => 9064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 8968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 753, 3 => 7326, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6291, 3 => 3833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2614, 3 => 7844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2303, 3 => 646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2075, 3 => 611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4687, 3 => 362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 8684, 3 => 9940, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4830, 3 => 2065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7038, 3 => 1363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1769, 3 => 7837, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3801, 3 => 1689, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10070, 3 => 2359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3667, 3 => 9918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1914, 3 => 6920, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4244, 3 => 5669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10245, 3 => 7821, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7648, 3 => 3944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3310, 3 => 5488, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6346, 3 => 9666, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7088, 3 => 6122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1291, 3 => 7827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 10592, 3 => 8945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3609, 3 => 7120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 9168, 3 => 9112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6203, 3 => 8052, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3330, 3 => 2895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4264, 3 => 10563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10556, 3 => 6496, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8807, 3 => 7645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1999, 3 => 4530, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9202, 3 => 6818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3403, 3 => 1734, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2106, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 24, 2 => 6881, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 25, 2 => 3895, 3 => 2171, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4062, 3 => 6424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 27, 2 => 3755, 3 => 9536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4683, 3 => 2131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7347, 3 => 8027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C8_9.csv, table is 160x46 (920.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9 : integer_2d_array_t(0 to 159)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 6235, 3 => 2848, 4 => 3222),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5800, 3 => 3492, 4 => 5348),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2757, 3 => 927, 4 => 90),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6961, 3 => 4516, 4 => 4739),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1172, 3 => 3237, 4 => 6264),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1927, 3 => 2425, 4 => 3683),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3714, 3 => 6309, 4 => 2495),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 3070, 3 => 6342, 4 => 7154),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2428, 3 => 613, 4 => 3761),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 2906, 3 => 264, 4 => 5927),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 1716, 3 => 1950, 4 => 4273),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4613, 3 => 6179, 4 => 3491),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 4865, 3 => 3286, 4 => 6005),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1343, 3 => 5923, 4 => 3529),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 4589, 3 => 4035, 4 => 2132),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 1579, 3 => 3920, 4 => 6737),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1644, 3 => 1191, 4 => 5998),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 1482, 3 => 2381, 4 => 4620),
    18 => integer_vector_t'(0 => 4, 1 => 18, 2 => 6791, 3 => 6014, 4 => 6596),
    19 => integer_vector_t'(0 => 4, 1 => 19, 2 => 2738, 3 => 5918, 4 => 3786),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5156, 3 => 6166, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1504, 3 => 4356, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 130, 3 => 1904, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6027, 3 => 3187, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6718, 3 => 759, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6240, 3 => 2870, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2343, 3 => 1311, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1039, 3 => 5465, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6617, 3 => 2513, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1588, 3 => 5222, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6561, 3 => 535, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4765, 3 => 2054, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5966, 3 => 6892, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1969, 3 => 3869, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3571, 3 => 2420, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4632, 3 => 981, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3215, 3 => 4163, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 17, 2 => 973, 3 => 3117, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 18, 2 => 3802, 3 => 6198, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3794, 3 => 3948, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3196, 3 => 6126, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 1, 2 => 573, 3 => 1909, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 2, 2 => 850, 3 => 4034, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5622, 3 => 1601, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6005, 3 => 524, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5251, 3 => 5783, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 6, 2 => 172, 3 => 2032, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1875, 3 => 2475, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 8, 2 => 497, 3 => 1291, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2566, 3 => 3430, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1249, 3 => 740, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2944, 3 => 1948, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6528, 3 => 2899, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2243, 3 => 3616, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 14, 2 => 867, 3 => 3733, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1374, 3 => 4702, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4698, 3 => 2285, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4760, 3 => 3917, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1859, 3 => 4058, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6141, 3 => 3527, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2148, 3 => 5066, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1306, 3 => 145, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2319, 3 => 871, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3463, 3 => 1061, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5554, 3 => 6647, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5837, 3 => 339, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5821, 3 => 4932, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6356, 3 => 4756, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3930, 3 => 418, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 211, 3 => 3094, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1007, 3 => 4928, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3584, 3 => 1235, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6982, 3 => 2869, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1612, 3 => 1013, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 953, 3 => 4964, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4555, 3 => 4410, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4925, 3 => 4842, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5778, 3 => 600, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6509, 3 => 2417, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1260, 3 => 4903, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3369, 3 => 3031, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3557, 3 => 3224, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3028, 3 => 583, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3258, 3 => 440, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6226, 3 => 6655, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4895, 3 => 1094, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1481, 3 => 6847, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4433, 3 => 1932, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2107, 3 => 1649, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2119, 3 => 2065, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4003, 3 => 6388, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6720, 3 => 3622, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3694, 3 => 4521, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1164, 3 => 7050, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1965, 3 => 3613, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4331, 3 => 66, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2970, 3 => 1796, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4652, 3 => 3218, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1762, 3 => 4777, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5736, 3 => 1399, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 0, 2 => 970, 3 => 2572, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2062, 3 => 6599, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4597, 3 => 4870, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1228, 3 => 6913, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4159, 3 => 1037, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2916, 3 => 2362, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 6, 2 => 395, 3 => 1226, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6911, 3 => 4548, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4618, 3 => 2241, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4120, 3 => 4280, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5825, 3 => 474, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2154, 3 => 5558, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3793, 3 => 5471, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5707, 3 => 1595, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1403, 3 => 325, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6601, 3 => 5183, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6369, 3 => 4569, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4846, 3 => 896, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 18, 2 => 7092, 3 => 6184, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6764, 3 => 7127, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6358, 3 => 1951, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3117, 3 => 6960, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2710, 3 => 7062, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1133, 3 => 3604, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3694, 3 => 657, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1355, 3 => 110, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3329, 3 => 6736, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2505, 3 => 3407, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2462, 3 => 4806, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4216, 3 => 214, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5348, 3 => 5619, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6627, 3 => 6243, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 2644, 3 => 5073, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4212, 3 => 5088, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3463, 3 => 3889, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5306, 3 => 478, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4320, 3 => 6121, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3961, 3 => 1125, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5699, 3 => 1195, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6511, 3 => 792, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3934, 3 => 2778, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3238, 3 => 6587, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1111, 3 => 6596, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1457, 3 => 6226, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1446, 3 => 3885, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3907, 3 => 4043, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6839, 3 => 2873, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1733, 3 => 5615, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5202, 3 => 4269, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3024, 3 => 4722, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5445, 3 => 6372, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 11, 2 => 370, 3 => 1828, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4695, 3 => 1600, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 13, 2 => 680, 3 => 2074, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1801, 3 => 6690, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2669, 3 => 1377, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2463, 3 => 1681, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5972, 3 => 5171, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5728, 3 => 4284, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1696, 3 => 1459, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C9_10.csv, table is 162x46 (931.5 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10 : integer_2d_array_t(0 to 161)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 5611, 3 => 2563, 4 => 2900),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5220, 3 => 3143, 4 => 4813),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2481, 3 => 834, 4 => 81),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6265, 3 => 4064, 4 => 4265),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1055, 3 => 2914, 4 => 5638),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1734, 3 => 2182, 4 => 3315),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3342, 3 => 5678, 4 => 2246),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 2185, 3 => 552, 4 => 3385),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2615, 3 => 236, 4 => 5334),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 1546, 3 => 1755, 4 => 3846),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 4154, 3 => 5561, 4 => 3142),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4382, 3 => 2957, 4 => 5400),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 1209, 3 => 5329, 4 => 3179),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1421, 3 => 3528, 4 => 6063),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 1480, 3 => 1072, 4 => 5398),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 3843, 3 => 1777, 4 => 4369),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1334, 3 => 2145, 4 => 4163),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 2368, 3 => 5055, 4 => 260),
    18 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6118, 3 => 5405, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2994, 3 => 4370, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3405, 3 => 1669, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4640, 3 => 5550, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1354, 3 => 3921, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 5, 2 => 117, 3 => 1713, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5425, 3 => 2866, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6047, 3 => 683, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5616, 3 => 2582, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2108, 3 => 1179, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 10, 2 => 933, 3 => 4921, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5953, 3 => 2261, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1430, 3 => 4699, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5905, 3 => 480, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4289, 3 => 1846, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5374, 3 => 6208, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1775, 3 => 3476, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3216, 3 => 2178, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4165, 3 => 884, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2896, 3 => 3744, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 2801, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3423, 3 => 5579, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3404, 3 => 3552, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2876, 3 => 5515, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 516, 3 => 1719, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 765, 3 => 3631, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5059, 3 => 1441, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5629, 3 => 598, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5405, 3 => 473, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4724, 3 => 5210, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 155, 3 => 1832, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1689, 3 => 2229, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 449, 3 => 1164, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2308, 3 => 3088, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1122, 3 => 669, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2268, 3 => 5758, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5878, 3 => 2609, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 1, 2 => 782, 3 => 3359, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1231, 3 => 4231, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4225, 3 => 2052, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4286, 3 => 3517, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5531, 3 => 3184, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1935, 3 => 4560, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1174, 3 => 131, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3115, 3 => 956, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3129, 3 => 1088, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5238, 3 => 4440, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5722, 3 => 4280, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3540, 3 => 375, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 13, 2 => 191, 3 => 2782, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 14, 2 => 906, 3 => 4432, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3225, 3 => 1111, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6296, 3 => 2583, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1457, 3 => 903, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 855, 3 => 4475, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4097, 3 => 3970, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4433, 3 => 4361, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5198, 3 => 541, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1146, 3 => 4426, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3202, 3 => 2902, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2724, 3 => 525, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1083, 3 => 4124, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2326, 3 => 6003, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5605, 3 => 5990, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4376, 3 => 1579, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4407, 3 => 984, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1332, 3 => 6163, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5359, 3 => 3975, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1907, 3 => 1854, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3601, 3 => 5748, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6056, 3 => 3266, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3322, 3 => 4085, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1768, 3 => 3244, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2149, 3 => 144, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1589, 3 => 4291, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5154, 3 => 1252, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1855, 3 => 5939, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4820, 3 => 2706, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1475, 3 => 3360, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4266, 3 => 693, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4156, 3 => 2018, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2103, 3 => 752, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3710, 3 => 3853, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5123, 3 => 931, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6146, 3 => 3323, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1939, 3 => 5002, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5140, 3 => 1437, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1263, 3 => 293, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5949, 3 => 4665, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4548, 3 => 6380, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3171, 3 => 4690, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5204, 3 => 2114, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6384, 3 => 5565, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5722, 3 => 1757, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2805, 3 => 6264, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1202, 3 => 2616, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1018, 3 => 3244, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4018, 3 => 5289, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2257, 3 => 3067, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2483, 3 => 3073, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1196, 3 => 5329, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 649, 3 => 3918, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3791, 3 => 4581, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5028, 3 => 3803, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3119, 3 => 3506, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4779, 3 => 431, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3888, 3 => 5510, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4387, 3 => 4084, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5836, 3 => 1692, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5126, 3 => 1078, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 2, 2 => 5721, 3 => 6165, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3540, 3 => 2499, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2225, 3 => 6348, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1044, 3 => 1484, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6323, 3 => 4042, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1313, 3 => 5603, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1303, 3 => 3496, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3516, 3 => 3639, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5161, 3 => 2293, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4682, 3 => 3845, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3045, 3 => 643, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2818, 3 => 2616, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3267, 3 => 649, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6236, 3 => 593, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 16, 2 => 646, 3 => 2948, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4213, 3 => 1442, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5779, 3 => 1596, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2403, 3 => 1237, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2217, 3 => 1514, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5609, 3 => 716, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5155, 3 => 3858, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1517, 3 => 1312, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2554, 3 => 3158, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5280, 3 => 2643, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4990, 3 => 1353, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5648, 3 => 1170, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1152, 3 => 4366, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3561, 3 => 5368, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3581, 3 => 1411, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5647, 3 => 4661, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1542, 3 => 5401, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5078, 3 => 2687, 4 => -1),
    160 => integer_vector_t'(0 => 3, 1 => 16, 2 => 316, 3 => 1755, 4 => -1),
    161 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3392, 3 => 1991, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_2.csv, table is 20x100 (250.0 bytes)
  -- Resource estimation: 6 x 18 kB BRAMs or 3 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 5, 2 => 14, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_2 : integer_2d_array_t(0 to 19)(0 to 8) := (
    0 => integer_vector_t'(0 => 8, 1 => 20, 2 => 712, 3 => 2386, 4 => 6354, 5 => 4061, 6 => 1062, 7 => 5045, 8 => 5158),
    1 => integer_vector_t'(0 => 8, 1 => 21, 2 => 2543, 3 => 5748, 4 => 4822, 5 => 2348, 6 => 3089, 7 => 6328, 8 => 5876),
    2 => integer_vector_t'(0 => 8, 1 => 22, 2 => 926, 3 => 5701, 4 => 269, 5 => 3693, 6 => 2438, 7 => 3190, 8 => 3507),
    3 => integer_vector_t'(0 => 8, 1 => 23, 2 => 2802, 3 => 4520, 4 => 3577, 5 => 5324, 6 => 1091, 7 => 4667, 8 => 4449),
    4 => integer_vector_t'(0 => 8, 1 => 24, 2 => 5140, 3 => 2003, 4 => 1263, 5 => 4742, 6 => 6497, 7 => 1185, 8 => 6202),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4046, 3 => 6934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2855, 3 => 66, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6694, 3 => 212, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3439, 3 => 1158, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3850, 3 => 4422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5924, 3 => 290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1467, 3 => 4049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7820, 3 => 2242, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4606, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4633, 3 => 7877, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3884, 3 => 6868, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8935, 3 => 4996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3028, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5988, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7411, 3 => 3450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_3.csv, table is 15x170 (318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 13, 9 => 14, 10 => 14, 11 => 14, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_3 : integer_2d_array_t(0 to 14)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 416, 2 => 8909, 3 => 4156, 4 => 3216, 5 => 3112, 6 => 2560, 7 => 2912, 8 => 6405, 9 => 8593, 10 => 4969, 11 => 6723, 12 => 6912),
    1 => integer_vector_t'(0 => 12, 1 => 8978, 2 => 3011, 3 => 4339, 4 => 9312, 5 => 6396, 6 => 2957, 7 => 7288, 8 => 5485, 9 => 6031, 10 => 10218, 11 => 2226, 12 => 3575),
    2 => integer_vector_t'(0 => 12, 1 => 3383, 2 => 10059, 3 => 1114, 4 => 10008, 5 => 10147, 6 => 9384, 7 => 4290, 8 => 434, 9 => 5139, 10 => 3536, 11 => 1965, 12 => 2291),
    3 => integer_vector_t'(0 => 12, 1 => 2797, 2 => 3693, 3 => 7615, 4 => 7077, 5 => 743, 6 => 1941, 7 => 8716, 8 => 6215, 9 => 3840, 10 => 5140, 11 => 4582, 12 => 5420),
    4 => integer_vector_t'(0 => 12, 1 => 6110, 2 => 8551, 3 => 1515, 4 => 7404, 5 => 4879, 6 => 4946, 7 => 5383, 8 => 1831, 9 => 3441, 10 => 9569, 11 => 10472, 12 => 4306),
    5 => integer_vector_t'(0 => 3, 1 => 1505, 2 => 5682, 3 => 7778, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 7172, 2 => 6830, 3 => 6623, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7281, 2 => 3941, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 10270, 2 => 8669, 3 => 914, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 3622, 2 => 7563, 3 => 9388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 9930, 2 => 5058, 3 => 4554, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 4844, 2 => 9609, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 6883, 2 => 3237, 3 => 1714, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4768, 2 => 3878, 3 => 10017, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 10127, 2 => 3334, 3 => 8267, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_4.csv, table is 9x171 (192.375 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 13, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_4 : integer_2d_array_t(0 to 8)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 6295, 2 => 9626, 3 => 304, 4 => 7695, 5 => 4839, 6 => 4936, 7 => 1660, 8 => 144, 9 => 11203, 10 => 5567, 11 => 6347, 12 => 12557),
    1 => integer_vector_t'(0 => 12, 1 => 10691, 2 => 4988, 3 => 3859, 4 => 3734, 5 => 3071, 6 => 3494, 7 => 7687, 8 => 10313, 9 => 5964, 10 => 8069, 11 => 8296, 12 => 11090),
    2 => integer_vector_t'(0 => 12, 1 => 10774, 2 => 3613, 3 => 5208, 4 => 11177, 5 => 7676, 6 => 3549, 7 => 8746, 8 => 6583, 9 => 7239, 10 => 12265, 11 => 2674, 12 => 4292),
    3 => integer_vector_t'(0 => 12, 1 => 11869, 2 => 3708, 3 => 5981, 4 => 8718, 5 => 4908, 6 => 10650, 7 => 6805, 8 => 3334, 9 => 2627, 10 => 10461, 11 => 9285, 12 => 11120),
    4 => integer_vector_t'(0 => 3, 1 => 7844, 2 => 3079, 3 => 10773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 3385, 2 => 10854, 3 => 5747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1360, 2 => 12010, 3 => 12202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 6189, 2 => 4241, 3 => 2343, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9840, 2 => 12726, 3 => 4977, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_3.csv, table is 30x156 (585.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 13, 4 => 12, 5 => 12, 6 => 11, 7 => 12, 8 => 13, 9 => 12, 10 => 13, 11 => 12, 12 => 13, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_3 : integer_2d_array_t(0 to 29)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 2084, 3 => 1613, 4 => 1548, 5 => 1286, 6 => 1460, 7 => 3196, 8 => 4297, 9 => 2481, 10 => 3369, 11 => 3451, 12 => 4620, 13 => 2622),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 122, 3 => 1516, 4 => 3448, 5 => 2880, 6 => 1407, 7 => 1847, 8 => 3799, 9 => 3529, 10 => 373, 11 => 971, 12 => 4358, 13 => 3108),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 259, 3 => 3399, 4 => 929, 5 => 2650, 6 => 864, 7 => 3996, 8 => 3833, 9 => 107, 10 => 5287, 11 => 164, 12 => 3125, 13 => 2350),
    3 => integer_vector_t'(0 => 3, 1 => 3, 2 => 342, 3 => 3529, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4198, 3 => 2147, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1880, 3 => 4836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3864, 3 => 4910, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7, 2 => 243, 3 => 1542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3011, 3 => 1436, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2167, 3 => 2512, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4606, 3 => 1003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2835, 3 => 705, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3426, 3 => 2365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3848, 3 => 2474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1360, 3 => 1743, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 163, 3 => 2536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2583, 3 => 1180, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1542, 3 => 509, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4418, 3 => 1005, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5212, 3 => 5117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2155, 3 => 2922, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 347, 3 => 2696, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 226, 3 => 4296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1560, 3 => 487, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3926, 3 => 1640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 10, 2 => 149, 3 => 2928, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2364, 3 => 563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 12, 2 => 635, 3 => 688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 13, 2 => 231, 3 => 1684, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1129, 3 => 3894, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_5.csv, table is 18x168 (378.0 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 13, 8 => 13, 9 => 13, 10 => 14, 11 => 13, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_5 : integer_2d_array_t(0 to 17)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 5650, 2 => 4143, 3 => 8750, 4 => 583, 5 => 6720, 6 => 8071, 7 => 635, 8 => 1767, 9 => 1344, 10 => 6922, 11 => 738, 12 => 6658),
    1 => integer_vector_t'(0 => 12, 1 => 5696, 2 => 1685, 3 => 3207, 4 => 415, 5 => 7019, 6 => 5023, 7 => 5608, 8 => 2605, 9 => 857, 10 => 6915, 11 => 1770, 12 => 8016),
    2 => integer_vector_t'(0 => 12, 1 => 3992, 2 => 771, 3 => 2190, 4 => 7258, 5 => 8970, 6 => 7792, 7 => 1802, 8 => 1866, 9 => 6137, 10 => 8841, 11 => 886, 12 => 1931),
    3 => integer_vector_t'(0 => 12, 1 => 4108, 2 => 3781, 3 => 7577, 4 => 6810, 5 => 9322, 6 => 8226, 7 => 5396, 8 => 5867, 9 => 4428, 10 => 8827, 11 => 7766, 12 => 2254),
    4 => integer_vector_t'(0 => 12, 1 => 4247, 2 => 888, 3 => 4367, 4 => 8821, 5 => 9660, 6 => 324, 7 => 5864, 8 => 4774, 9 => 227, 10 => 7889, 11 => 6405, 12 => 8963),
    5 => integer_vector_t'(0 => 12, 1 => 9693, 2 => 500, 3 => 2520, 4 => 2227, 5 => 1811, 6 => 9330, 7 => 1928, 8 => 5140, 9 => 4030, 10 => 4824, 11 => 806, 12 => 3134),
    6 => integer_vector_t'(0 => 3, 1 => 1652, 2 => 8171, 3 => 1435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 3366, 2 => 6543, 3 => 3745, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9286, 2 => 8509, 3 => 4645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 7397, 2 => 5790, 3 => 8972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 6597, 2 => 4422, 3 => 1799, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 9276, 2 => 4041, 3 => 3847, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 8683, 2 => 7378, 3 => 4946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 5348, 2 => 1993, 3 => 9186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 6724, 2 => 9015, 3 => 5646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 4502, 2 => 4439, 3 => 8474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 5107, 2 => 7342, 3 => 9442, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 1387, 2 => 8910, 3 => 2660, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_4.csv, table is 33x133 (548.625 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 12, 4 => 13, 5 => 11, 6 => 10, 7 => 12, 8 => 11, 9 => 12, 10 => 10, 11 => 10, 12 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_4 : integer_2d_array_t(0 to 32)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 3, 2 => 3198, 3 => 478, 4 => 4207, 5 => 1481, 6 => 1009, 7 => 2616, 8 => 1924, 9 => 3437, 10 => 554, 11 => 683, 12 => 1801),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2681, 3 => 2135, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3107, 3 => 4027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2637, 3 => 3373, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 3830, 3 => 3449, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4129, 3 => 2060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4184, 3 => 2742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3946, 3 => 1070, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2239, 3 => 984, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1458, 3 => 3031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3003, 3 => 1328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1137, 3 => 1716, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 132, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1817, 3 => 638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1774, 3 => 3447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3632, 3 => 1257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 542, 3 => 3694, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1015, 3 => 1945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1948, 3 => 412, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 995, 3 => 2238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4141, 3 => 1907, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2480, 3 => 3079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3021, 3 => 1088, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 713, 3 => 1379, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 997, 3 => 3903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2323, 3 => 3361, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1110, 3 => 986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2532, 3 => 142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1690, 3 => 2405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1298, 3 => 1881, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 9, 2 => 615, 3 => 174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1648, 3 => 3112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1415, 3 => 2808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_5.csv, table is 27x160 (540.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 13, 2 => 13, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13, 9 => 13, 10 => 13, 11 => 13, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_5 : integer_2d_array_t(0 to 26)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 2765, 2 => 5713, 3 => 6426, 4 => 3596, 5 => 1374, 6 => 4811, 7 => 2182, 8 => 544, 9 => 3394, 10 => 2840, 11 => 4310, 12 => 771),
    1 => integer_vector_t'(0 => 12, 1 => 4951, 2 => 211, 3 => 2208, 4 => 723, 5 => 1246, 6 => 2928, 7 => 398, 8 => 5739, 9 => 265, 10 => 5601, 11 => 5993, 12 => 2615),
    2 => integer_vector_t'(0 => 12, 1 => 210, 2 => 4730, 3 => 5777, 4 => 3096, 5 => 4282, 6 => 6238, 7 => 4939, 8 => 1119, 9 => 6463, 10 => 5298, 11 => 6320, 12 => 4016),
    3 => integer_vector_t'(0 => 12, 1 => 4167, 2 => 2063, 3 => 4757, 4 => 3157, 5 => 5664, 6 => 3956, 7 => 6045, 8 => 563, 9 => 4284, 10 => 2441, 11 => 3412, 12 => 6334),
    4 => integer_vector_t'(0 => 12, 1 => 4201, 2 => 2428, 3 => 4474, 4 => 59, 5 => 1721, 6 => 736, 7 => 2997, 8 => 428, 9 => 3807, 10 => 1513, 11 => 4732, 12 => 6195),
    5 => integer_vector_t'(0 => 12, 1 => 2670, 2 => 3081, 3 => 5139, 4 => 3736, 5 => 1999, 6 => 5889, 7 => 4362, 8 => 3806, 9 => 4534, 10 => 5409, 11 => 6384, 12 => 5809),
    6 => integer_vector_t'(0 => 12, 1 => 5516, 2 => 1622, 3 => 2906, 4 => 3285, 5 => 1257, 6 => 5797, 7 => 3816, 8 => 817, 9 => 875, 10 => 2311, 11 => 3543, 12 => 1205),
    7 => integer_vector_t'(0 => 12, 1 => 4244, 2 => 2184, 3 => 5415, 4 => 1705, 5 => 5642, 6 => 4886, 7 => 2333, 8 => 287, 9 => 1848, 10 => 1121, 11 => 3595, 12 => 6022),
    8 => integer_vector_t'(0 => 12, 1 => 2142, 2 => 2830, 3 => 4069, 4 => 5654, 5 => 1295, 6 => 2951, 7 => 3919, 8 => 1356, 9 => 884, 10 => 1786, 11 => 396, 12 => 4738),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2161, 3 => 2653, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1380, 3 => 1461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2502, 3 => 3707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3971, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5985, 3 => 6062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1733, 3 => 6028, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3786, 3 => 1936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4292, 3 => 956, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5692, 3 => 3417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 266, 3 => 4878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4913, 3 => 3247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4763, 3 => 3937, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3590, 3 => 2903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2566, 3 => 4215, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5208, 3 => 4707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3940, 3 => 3388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5109, 3 => 4556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4908, 3 => 4177, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C4_5.csv, table is 35x30 (131.25 bytes)
  -- Resource estimation: 2 x 18 kB BRAMs or 1 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 4, 2 => 12, 3 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C4_5 : integer_2d_array_t(0 to 34)(0 to 3) := (
    0 => integer_vector_t'(0 => 3, 1 => 5, 2 => 896, 3 => 1565),
    1 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2493, 3 => 184),
    2 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 3210),
    3 => integer_vector_t'(0 => 3, 1 => 8, 2 => 727, 3 => 1339),
    4 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3428, 3 => 612),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2663, 3 => 1947),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 230, 3 => 2695),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2025, 3 => 2794),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3039, 3 => 283),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 862, 3 => 2889),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 376, 3 => 2110),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2034, 3 => 2286),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 951, 3 => 2068),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3108, 3 => 3542),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 307, 3 => 1421),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2272, 3 => 1197),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1800, 3 => 3280),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 331, 3 => 2308),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 465, 3 => 2552),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1038, 3 => 2479),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1383, 3 => 343),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 94, 3 => 236),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2619, 3 => 121),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1497, 3 => 2774),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2116, 3 => 1855),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 722, 3 => 1584),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2767, 3 => 1881),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2701, 3 => 1610),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3283, 3 => 1732),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 168, 3 => 1099),
    30 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3074, 3 => 243),
    31 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3460, 3 => 945),
    32 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2049, 3 => 1746),
    33 => integer_vector_t'(0 => 3, 1 => 8, 2 => 566, 3 => 1427),
    34 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3545, 3 => 1168)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C5_6.csv, table is 37x139 (642.875 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 3, 2 => 12, 3 => 12, 4 => 11, 5 => 10, 6 => 10, 7 => 10, 8 => 11, 9 => 9, 10 => 12, 11 => 12, 12 => 11, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C5_6 : integer_2d_array_t(0 to 36)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 3, 2 => 2409, 3 => 499, 4 => 1481, 5 => 908, 6 => 559, 7 => 716, 8 => 1270, 9 => 333, 10 => 2508, 11 => 2264, 12 => 1702, 13 => 2805),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2447, 3 => 1926, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 414, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2114, 3 => 842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 573, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2383, 3 => 2112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2286, 3 => 2348, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 545, 3 => 819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1264, 3 => 143, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1701, 3 => 2258, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 964, 3 => 166, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 114, 3 => 2413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2243, 3 => 81, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1245, 3 => 1581, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 1, 2 => 775, 3 => 169, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1696, 3 => 1104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1914, 3 => 2831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 4, 2 => 532, 3 => 1450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 5, 2 => 91, 3 => 974, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 6, 2 => 497, 3 => 2228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2326, 3 => 1579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2482, 3 => 256, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1117, 3 => 1261, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1257, 3 => 1658, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1478, 3 => 1225, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2511, 3 => 980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2320, 3 => 2675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 435, 3 => 1278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 228, 3 => 503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1885, 3 => 2369, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 1, 2 => 57, 3 => 483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 2, 2 => 838, 3 => 1050, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1231, 3 => 1990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1738, 3 => 68, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2392, 3 => 951, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 6, 2 => 163, 3 => 645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2644, 3 => 1704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C8_9.csv, table is 40x37 (185.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 2, 2 => 11, 3 => 11, 4 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C8_9 : integer_2d_array_t(0 to 39)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 1558, 3 => 712, 4 => 805),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 1450, 3 => 873, 4 => 1337),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 1741, 3 => 1129, 4 => 1184),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 294, 3 => 806, 4 => 1566),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 482, 3 => 605, 4 => 923),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 926, 3 => 1578, 4 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 777, 3 => 1374, 4 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 608, 3 => 151, 4 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1195, 3 => 210, 4 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1484, 3 => 692, 4 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 0, 2 => 427, 3 => 488, 4 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 1, 2 => 828, 3 => 1124, 4 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 1366, 4 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1500, 3 => 835, 4 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1496, 3 => 502, 4 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1006, 3 => 1701, 4 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1155, 3 => 97, 4 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 657, 3 => 1403, 4 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1453, 3 => 624, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 429, 3 => 1495, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 809, 3 => 385, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 367, 3 => 151, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1323, 3 => 202, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 960, 3 => 318, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1451, 3 => 1039, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1098, 3 => 1722, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1015, 3 => 1428, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1261, 3 => 1564, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 544, 3 => 1190, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1472, 3 => 1246, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 508, 3 => 630, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 421, 3 => 1704, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 284, 3 => 898, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 392, 3 => 577, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1155, 3 => 556, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 0, 2 => 631, 3 => 1000, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 1, 2 => 732, 3 => 1368, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1328, 3 => 329, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1515, 3 => 506, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1104, 3 => 1172, 4 => -1)
  );


  -- Record with LDPC metadata
  type ldpc_metadata_t is record
    addr : integer;
    q : integer;
    stage_0_loops: integer;
    stage_0_rows: integer;
    stage_1_loops: integer;
    stage_1_rows: integer;
  end record ldpc_metadata_t;

  -- Reduce the footprint of this
  constant LDPC_TABLE_DATA_WIDTH : integer := numbits(max(DVB_N_LDPC));

  -- Use this function to get the starting address of a given config within the LDPC_DATA_TABLE
  function get_ldpc_metadata (
    constant frame_length : frame_type_t;
    constant code_rate : code_rate_t) return ldpc_metadata_t;


  constant LDPC_DATA_TABLE : std_logic_vector_2d_t(0 to 6446)(16 - 1 downto 0) := (
    -- Table for fecframe_normal, C1_2
       0 => std_logic_vector(to_unsigned(   54, 16)), --    54 / 0x0036
       1 => std_logic_vector(to_unsigned( 9318, 16)), --  9318 / 0x2466
       2 => std_logic_vector(to_unsigned(14392, 16)), -- 14392 / 0x3838
       3 => std_logic_vector(to_unsigned(27561, 16)), -- 27561 / 0x6ba9
       4 => std_logic_vector(to_unsigned(26909, 16)), -- 26909 / 0x691d
       5 => std_logic_vector(to_unsigned(10219, 16)), -- 10219 / 0x27eb
       6 => std_logic_vector(to_unsigned( 2534, 16)), --  2534 / 0x09e6
       7 => std_logic_vector(to_unsigned( 8597, 16)), --  8597 / 0x2195 -- last item of row
       8 => std_logic_vector(to_unsigned(   55, 16)), --    55 / 0x0037
       9 => std_logic_vector(to_unsigned( 7263, 16)), --  7263 / 0x1c5f
      10 => std_logic_vector(to_unsigned( 4635, 16)), --  4635 / 0x121b
      11 => std_logic_vector(to_unsigned( 2530, 16)), --  2530 / 0x09e2
      12 => std_logic_vector(to_unsigned(28130, 16)), -- 28130 / 0x6de2
      13 => std_logic_vector(to_unsigned( 3033, 16)), --  3033 / 0x0bd9
      14 => std_logic_vector(to_unsigned(23830, 16)), -- 23830 / 0x5d16
      15 => std_logic_vector(to_unsigned( 3651, 16)), --  3651 / 0x0e43 -- last item of row
      16 => std_logic_vector(to_unsigned(   56, 16)), --    56 / 0x0038
      17 => std_logic_vector(to_unsigned(24731, 16)), -- 24731 / 0x609b
      18 => std_logic_vector(to_unsigned(23583, 16)), -- 23583 / 0x5c1f
      19 => std_logic_vector(to_unsigned(26036, 16)), -- 26036 / 0x65b4
      20 => std_logic_vector(to_unsigned(17299, 16)), -- 17299 / 0x4393
      21 => std_logic_vector(to_unsigned( 5750, 16)), --  5750 / 0x1676
      22 => std_logic_vector(to_unsigned(  792, 16)), --   792 / 0x0318
      23 => std_logic_vector(to_unsigned( 9169, 16)), --  9169 / 0x23d1 -- last item of row
      24 => std_logic_vector(to_unsigned(   57, 16)), --    57 / 0x0039
      25 => std_logic_vector(to_unsigned( 5811, 16)), --  5811 / 0x16b3
      26 => std_logic_vector(to_unsigned(26154, 16)), -- 26154 / 0x662a
      27 => std_logic_vector(to_unsigned(18653, 16)), -- 18653 / 0x48dd
      28 => std_logic_vector(to_unsigned(11551, 16)), -- 11551 / 0x2d1f
      29 => std_logic_vector(to_unsigned(15447, 16)), -- 15447 / 0x3c57
      30 => std_logic_vector(to_unsigned(13685, 16)), -- 13685 / 0x3575
      31 => std_logic_vector(to_unsigned(16264, 16)), -- 16264 / 0x3f88 -- last item of row
      32 => std_logic_vector(to_unsigned(   58, 16)), --    58 / 0x003a
      33 => std_logic_vector(to_unsigned(12610, 16)), -- 12610 / 0x3142
      34 => std_logic_vector(to_unsigned(11347, 16)), -- 11347 / 0x2c53
      35 => std_logic_vector(to_unsigned(28768, 16)), -- 28768 / 0x7060
      36 => std_logic_vector(to_unsigned( 2792, 16)), --  2792 / 0x0ae8
      37 => std_logic_vector(to_unsigned( 3174, 16)), --  3174 / 0x0c66
      38 => std_logic_vector(to_unsigned(29371, 16)), -- 29371 / 0x72bb
      39 => std_logic_vector(to_unsigned(12997, 16)), -- 12997 / 0x32c5 -- last item of row
      40 => std_logic_vector(to_unsigned(   59, 16)), --    59 / 0x003b
      41 => std_logic_vector(to_unsigned(16789, 16)), -- 16789 / 0x4195
      42 => std_logic_vector(to_unsigned(16018, 16)), -- 16018 / 0x3e92
      43 => std_logic_vector(to_unsigned(21449, 16)), -- 21449 / 0x53c9
      44 => std_logic_vector(to_unsigned( 6165, 16)), --  6165 / 0x1815
      45 => std_logic_vector(to_unsigned(21202, 16)), -- 21202 / 0x52d2
      46 => std_logic_vector(to_unsigned(15850, 16)), -- 15850 / 0x3dea
      47 => std_logic_vector(to_unsigned( 3186, 16)), --  3186 / 0x0c72 -- last item of row
      48 => std_logic_vector(to_unsigned(   60, 16)), --    60 / 0x003c
      49 => std_logic_vector(to_unsigned(31016, 16)), -- 31016 / 0x7928
      50 => std_logic_vector(to_unsigned(21449, 16)), -- 21449 / 0x53c9
      51 => std_logic_vector(to_unsigned(17618, 16)), -- 17618 / 0x44d2
      52 => std_logic_vector(to_unsigned( 6213, 16)), --  6213 / 0x1845
      53 => std_logic_vector(to_unsigned(12166, 16)), -- 12166 / 0x2f86
      54 => std_logic_vector(to_unsigned( 8334, 16)), --  8334 / 0x208e
      55 => std_logic_vector(to_unsigned(18212, 16)), -- 18212 / 0x4724 -- last item of row
      56 => std_logic_vector(to_unsigned(   61, 16)), --    61 / 0x003d
      57 => std_logic_vector(to_unsigned(22836, 16)), -- 22836 / 0x5934
      58 => std_logic_vector(to_unsigned(14213, 16)), -- 14213 / 0x3785
      59 => std_logic_vector(to_unsigned(11327, 16)), -- 11327 / 0x2c3f
      60 => std_logic_vector(to_unsigned( 5896, 16)), --  5896 / 0x1708
      61 => std_logic_vector(to_unsigned(  718, 16)), --   718 / 0x02ce
      62 => std_logic_vector(to_unsigned(11727, 16)), -- 11727 / 0x2dcf
      63 => std_logic_vector(to_unsigned( 9308, 16)), --  9308 / 0x245c -- last item of row
      64 => std_logic_vector(to_unsigned(   62, 16)), --    62 / 0x003e
      65 => std_logic_vector(to_unsigned( 2091, 16)), --  2091 / 0x082b
      66 => std_logic_vector(to_unsigned(24941, 16)), -- 24941 / 0x616d
      67 => std_logic_vector(to_unsigned(29966, 16)), -- 29966 / 0x750e
      68 => std_logic_vector(to_unsigned(23634, 16)), -- 23634 / 0x5c52
      69 => std_logic_vector(to_unsigned( 9013, 16)), --  9013 / 0x2335
      70 => std_logic_vector(to_unsigned(15587, 16)), -- 15587 / 0x3ce3
      71 => std_logic_vector(to_unsigned( 5444, 16)), --  5444 / 0x1544 -- last item of row
      72 => std_logic_vector(to_unsigned(   63, 16)), --    63 / 0x003f
      73 => std_logic_vector(to_unsigned(22207, 16)), -- 22207 / 0x56bf
      74 => std_logic_vector(to_unsigned( 3983, 16)), --  3983 / 0x0f8f
      75 => std_logic_vector(to_unsigned(16904, 16)), -- 16904 / 0x4208
      76 => std_logic_vector(to_unsigned(28534, 16)), -- 28534 / 0x6f76
      77 => std_logic_vector(to_unsigned(21415, 16)), -- 21415 / 0x53a7
      78 => std_logic_vector(to_unsigned(27524, 16)), -- 27524 / 0x6b84
      79 => std_logic_vector(to_unsigned(25912, 16)), -- 25912 / 0x6538 -- last item of row
      80 => std_logic_vector(to_unsigned(   64, 16)), --    64 / 0x0040
      81 => std_logic_vector(to_unsigned(25687, 16)), -- 25687 / 0x6457
      82 => std_logic_vector(to_unsigned( 4501, 16)), --  4501 / 0x1195
      83 => std_logic_vector(to_unsigned(22193, 16)), -- 22193 / 0x56b1
      84 => std_logic_vector(to_unsigned(14665, 16)), -- 14665 / 0x3949
      85 => std_logic_vector(to_unsigned(14798, 16)), -- 14798 / 0x39ce
      86 => std_logic_vector(to_unsigned(16158, 16)), -- 16158 / 0x3f1e
      87 => std_logic_vector(to_unsigned( 5491, 16)), --  5491 / 0x1573 -- last item of row
      88 => std_logic_vector(to_unsigned(   65, 16)), --    65 / 0x0041
      89 => std_logic_vector(to_unsigned( 4520, 16)), --  4520 / 0x11a8
      90 => std_logic_vector(to_unsigned(17094, 16)), -- 17094 / 0x42c6
      91 => std_logic_vector(to_unsigned(23397, 16)), -- 23397 / 0x5b65
      92 => std_logic_vector(to_unsigned( 4264, 16)), --  4264 / 0x10a8
      93 => std_logic_vector(to_unsigned(22370, 16)), -- 22370 / 0x5762
      94 => std_logic_vector(to_unsigned(16941, 16)), -- 16941 / 0x422d
      95 => std_logic_vector(to_unsigned(21526, 16)), -- 21526 / 0x5416 -- last item of row
      96 => std_logic_vector(to_unsigned(   66, 16)), --    66 / 0x0042
      97 => std_logic_vector(to_unsigned(10490, 16)), -- 10490 / 0x28fa
      98 => std_logic_vector(to_unsigned( 6182, 16)), --  6182 / 0x1826
      99 => std_logic_vector(to_unsigned(32370, 16)), -- 32370 / 0x7e72
     100 => std_logic_vector(to_unsigned( 9597, 16)), --  9597 / 0x257d
     101 => std_logic_vector(to_unsigned(30841, 16)), -- 30841 / 0x7879
     102 => std_logic_vector(to_unsigned(25954, 16)), -- 25954 / 0x6562
     103 => std_logic_vector(to_unsigned( 2762, 16)), --  2762 / 0x0aca -- last item of row
     104 => std_logic_vector(to_unsigned(   67, 16)), --    67 / 0x0043
     105 => std_logic_vector(to_unsigned(22120, 16)), -- 22120 / 0x5668
     106 => std_logic_vector(to_unsigned(22865, 16)), -- 22865 / 0x5951
     107 => std_logic_vector(to_unsigned(29870, 16)), -- 29870 / 0x74ae
     108 => std_logic_vector(to_unsigned(15147, 16)), -- 15147 / 0x3b2b
     109 => std_logic_vector(to_unsigned(13668, 16)), -- 13668 / 0x3564
     110 => std_logic_vector(to_unsigned(14955, 16)), -- 14955 / 0x3a6b
     111 => std_logic_vector(to_unsigned(19235, 16)), -- 19235 / 0x4b23 -- last item of row
     112 => std_logic_vector(to_unsigned(   68, 16)), --    68 / 0x0044
     113 => std_logic_vector(to_unsigned( 6689, 16)), --  6689 / 0x1a21
     114 => std_logic_vector(to_unsigned(18408, 16)), -- 18408 / 0x47e8
     115 => std_logic_vector(to_unsigned(18346, 16)), -- 18346 / 0x47aa
     116 => std_logic_vector(to_unsigned( 9918, 16)), --  9918 / 0x26be
     117 => std_logic_vector(to_unsigned(25746, 16)), -- 25746 / 0x6492
     118 => std_logic_vector(to_unsigned( 5443, 16)), --  5443 / 0x1543
     119 => std_logic_vector(to_unsigned(20645, 16)), -- 20645 / 0x50a5 -- last item of row
     120 => std_logic_vector(to_unsigned(   69, 16)), --    69 / 0x0045
     121 => std_logic_vector(to_unsigned(29982, 16)), -- 29982 / 0x751e
     122 => std_logic_vector(to_unsigned(12529, 16)), -- 12529 / 0x30f1
     123 => std_logic_vector(to_unsigned(13858, 16)), -- 13858 / 0x3622
     124 => std_logic_vector(to_unsigned( 4746, 16)), --  4746 / 0x128a
     125 => std_logic_vector(to_unsigned(30370, 16)), -- 30370 / 0x76a2
     126 => std_logic_vector(to_unsigned(10023, 16)), -- 10023 / 0x2727
     127 => std_logic_vector(to_unsigned(24828, 16)), -- 24828 / 0x60fc -- last item of row
     128 => std_logic_vector(to_unsigned(   70, 16)), --    70 / 0x0046
     129 => std_logic_vector(to_unsigned( 1262, 16)), --  1262 / 0x04ee
     130 => std_logic_vector(to_unsigned(28032, 16)), -- 28032 / 0x6d80
     131 => std_logic_vector(to_unsigned(29888, 16)), -- 29888 / 0x74c0
     132 => std_logic_vector(to_unsigned(13063, 16)), -- 13063 / 0x3307
     133 => std_logic_vector(to_unsigned(24033, 16)), -- 24033 / 0x5de1
     134 => std_logic_vector(to_unsigned(21951, 16)), -- 21951 / 0x55bf
     135 => std_logic_vector(to_unsigned( 7863, 16)), --  7863 / 0x1eb7 -- last item of row
     136 => std_logic_vector(to_unsigned(   71, 16)), --    71 / 0x0047
     137 => std_logic_vector(to_unsigned( 6594, 16)), --  6594 / 0x19c2
     138 => std_logic_vector(to_unsigned(29642, 16)), -- 29642 / 0x73ca
     139 => std_logic_vector(to_unsigned(31451, 16)), -- 31451 / 0x7adb
     140 => std_logic_vector(to_unsigned(14831, 16)), -- 14831 / 0x39ef
     141 => std_logic_vector(to_unsigned( 9509, 16)), --  9509 / 0x2525
     142 => std_logic_vector(to_unsigned( 9335, 16)), --  9335 / 0x2477
     143 => std_logic_vector(to_unsigned(31552, 16)), -- 31552 / 0x7b40 -- last item of row
     144 => std_logic_vector(to_unsigned(   72, 16)), --    72 / 0x0048
     145 => std_logic_vector(to_unsigned( 1358, 16)), --  1358 / 0x054e
     146 => std_logic_vector(to_unsigned( 6454, 16)), --  6454 / 0x1936
     147 => std_logic_vector(to_unsigned(16633, 16)), -- 16633 / 0x40f9
     148 => std_logic_vector(to_unsigned(20354, 16)), -- 20354 / 0x4f82
     149 => std_logic_vector(to_unsigned(24598, 16)), -- 24598 / 0x6016
     150 => std_logic_vector(to_unsigned(  624, 16)), --   624 / 0x0270
     151 => std_logic_vector(to_unsigned( 5265, 16)), --  5265 / 0x1491 -- last item of row
     152 => std_logic_vector(to_unsigned(   73, 16)), --    73 / 0x0049
     153 => std_logic_vector(to_unsigned(19529, 16)), -- 19529 / 0x4c49
     154 => std_logic_vector(to_unsigned(  295, 16)), --   295 / 0x0127
     155 => std_logic_vector(to_unsigned(18011, 16)), -- 18011 / 0x465b
     156 => std_logic_vector(to_unsigned( 3080, 16)), --  3080 / 0x0c08
     157 => std_logic_vector(to_unsigned(13364, 16)), -- 13364 / 0x3434
     158 => std_logic_vector(to_unsigned( 8032, 16)), --  8032 / 0x1f60
     159 => std_logic_vector(to_unsigned(15323, 16)), -- 15323 / 0x3bdb -- last item of row
     160 => std_logic_vector(to_unsigned(   74, 16)), --    74 / 0x004a
     161 => std_logic_vector(to_unsigned(11981, 16)), -- 11981 / 0x2ecd
     162 => std_logic_vector(to_unsigned( 1510, 16)), --  1510 / 0x05e6
     163 => std_logic_vector(to_unsigned( 7960, 16)), --  7960 / 0x1f18
     164 => std_logic_vector(to_unsigned(21462, 16)), -- 21462 / 0x53d6
     165 => std_logic_vector(to_unsigned( 9129, 16)), --  9129 / 0x23a9
     166 => std_logic_vector(to_unsigned(11370, 16)), -- 11370 / 0x2c6a
     167 => std_logic_vector(to_unsigned(25741, 16)), -- 25741 / 0x648d -- last item of row
     168 => std_logic_vector(to_unsigned(   75, 16)), --    75 / 0x004b
     169 => std_logic_vector(to_unsigned( 9276, 16)), --  9276 / 0x243c
     170 => std_logic_vector(to_unsigned(29656, 16)), -- 29656 / 0x73d8
     171 => std_logic_vector(to_unsigned( 4543, 16)), --  4543 / 0x11bf
     172 => std_logic_vector(to_unsigned(30699, 16)), -- 30699 / 0x77eb
     173 => std_logic_vector(to_unsigned(20646, 16)), -- 20646 / 0x50a6
     174 => std_logic_vector(to_unsigned(21921, 16)), -- 21921 / 0x55a1
     175 => std_logic_vector(to_unsigned(28050, 16)), -- 28050 / 0x6d92 -- last item of row
     176 => std_logic_vector(to_unsigned(   76, 16)), --    76 / 0x004c
     177 => std_logic_vector(to_unsigned(15975, 16)), -- 15975 / 0x3e67
     178 => std_logic_vector(to_unsigned(25634, 16)), -- 25634 / 0x6422
     179 => std_logic_vector(to_unsigned( 5520, 16)), --  5520 / 0x1590
     180 => std_logic_vector(to_unsigned(31119, 16)), -- 31119 / 0x798f
     181 => std_logic_vector(to_unsigned(13715, 16)), -- 13715 / 0x3593
     182 => std_logic_vector(to_unsigned(21949, 16)), -- 21949 / 0x55bd
     183 => std_logic_vector(to_unsigned(19605, 16)), -- 19605 / 0x4c95 -- last item of row
     184 => std_logic_vector(to_unsigned(   77, 16)), --    77 / 0x004d
     185 => std_logic_vector(to_unsigned(18688, 16)), -- 18688 / 0x4900
     186 => std_logic_vector(to_unsigned( 4608, 16)), --  4608 / 0x1200
     187 => std_logic_vector(to_unsigned(31755, 16)), -- 31755 / 0x7c0b
     188 => std_logic_vector(to_unsigned(30165, 16)), -- 30165 / 0x75d5
     189 => std_logic_vector(to_unsigned(13103, 16)), -- 13103 / 0x332f
     190 => std_logic_vector(to_unsigned(10706, 16)), -- 10706 / 0x29d2
     191 => std_logic_vector(to_unsigned(29224, 16)), -- 29224 / 0x7228 -- last item of row
     192 => std_logic_vector(to_unsigned(   78, 16)), --    78 / 0x004e
     193 => std_logic_vector(to_unsigned(21514, 16)), -- 21514 / 0x540a
     194 => std_logic_vector(to_unsigned(23117, 16)), -- 23117 / 0x5a4d
     195 => std_logic_vector(to_unsigned(12245, 16)), -- 12245 / 0x2fd5
     196 => std_logic_vector(to_unsigned(26035, 16)), -- 26035 / 0x65b3
     197 => std_logic_vector(to_unsigned(31656, 16)), -- 31656 / 0x7ba8
     198 => std_logic_vector(to_unsigned(25631, 16)), -- 25631 / 0x641f
     199 => std_logic_vector(to_unsigned(30699, 16)), -- 30699 / 0x77eb -- last item of row
     200 => std_logic_vector(to_unsigned(   79, 16)), --    79 / 0x004f
     201 => std_logic_vector(to_unsigned( 9674, 16)), --  9674 / 0x25ca
     202 => std_logic_vector(to_unsigned(24966, 16)), -- 24966 / 0x6186
     203 => std_logic_vector(to_unsigned(31285, 16)), -- 31285 / 0x7a35
     204 => std_logic_vector(to_unsigned(29908, 16)), -- 29908 / 0x74d4
     205 => std_logic_vector(to_unsigned(17042, 16)), -- 17042 / 0x4292
     206 => std_logic_vector(to_unsigned(24588, 16)), -- 24588 / 0x600c
     207 => std_logic_vector(to_unsigned(31857, 16)), -- 31857 / 0x7c71 -- last item of row
     208 => std_logic_vector(to_unsigned(   80, 16)), --    80 / 0x0050
     209 => std_logic_vector(to_unsigned(21856, 16)), -- 21856 / 0x5560
     210 => std_logic_vector(to_unsigned(27777, 16)), -- 27777 / 0x6c81
     211 => std_logic_vector(to_unsigned(29919, 16)), -- 29919 / 0x74df
     212 => std_logic_vector(to_unsigned(27000, 16)), -- 27000 / 0x6978
     213 => std_logic_vector(to_unsigned(14897, 16)), -- 14897 / 0x3a31
     214 => std_logic_vector(to_unsigned(11409, 16)), -- 11409 / 0x2c91
     215 => std_logic_vector(to_unsigned( 7122, 16)), --  7122 / 0x1bd2 -- last item of row
     216 => std_logic_vector(to_unsigned(   81, 16)), --    81 / 0x0051
     217 => std_logic_vector(to_unsigned(29773, 16)), -- 29773 / 0x744d
     218 => std_logic_vector(to_unsigned(23310, 16)), -- 23310 / 0x5b0e
     219 => std_logic_vector(to_unsigned(  263, 16)), --   263 / 0x0107
     220 => std_logic_vector(to_unsigned( 4877, 16)), --  4877 / 0x130d
     221 => std_logic_vector(to_unsigned(28622, 16)), -- 28622 / 0x6fce
     222 => std_logic_vector(to_unsigned(20545, 16)), -- 20545 / 0x5041
     223 => std_logic_vector(to_unsigned(22092, 16)), -- 22092 / 0x564c -- last item of row
     224 => std_logic_vector(to_unsigned(   82, 16)), --    82 / 0x0052
     225 => std_logic_vector(to_unsigned(15605, 16)), -- 15605 / 0x3cf5
     226 => std_logic_vector(to_unsigned( 5651, 16)), --  5651 / 0x1613
     227 => std_logic_vector(to_unsigned(21864, 16)), -- 21864 / 0x5568
     228 => std_logic_vector(to_unsigned( 3967, 16)), --  3967 / 0x0f7f
     229 => std_logic_vector(to_unsigned(14419, 16)), -- 14419 / 0x3853
     230 => std_logic_vector(to_unsigned(22757, 16)), -- 22757 / 0x58e5
     231 => std_logic_vector(to_unsigned(15896, 16)), -- 15896 / 0x3e18 -- last item of row
     232 => std_logic_vector(to_unsigned(   83, 16)), --    83 / 0x0053
     233 => std_logic_vector(to_unsigned(30145, 16)), -- 30145 / 0x75c1
     234 => std_logic_vector(to_unsigned( 1759, 16)), --  1759 / 0x06df
     235 => std_logic_vector(to_unsigned(10139, 16)), -- 10139 / 0x279b
     236 => std_logic_vector(to_unsigned(29223, 16)), -- 29223 / 0x7227
     237 => std_logic_vector(to_unsigned(26086, 16)), -- 26086 / 0x65e6
     238 => std_logic_vector(to_unsigned(10556, 16)), -- 10556 / 0x293c
     239 => std_logic_vector(to_unsigned( 5098, 16)), --  5098 / 0x13ea -- last item of row
     240 => std_logic_vector(to_unsigned(   84, 16)), --    84 / 0x0054
     241 => std_logic_vector(to_unsigned(18815, 16)), -- 18815 / 0x497f
     242 => std_logic_vector(to_unsigned(16575, 16)), -- 16575 / 0x40bf
     243 => std_logic_vector(to_unsigned( 2936, 16)), --  2936 / 0x0b78
     244 => std_logic_vector(to_unsigned(24457, 16)), -- 24457 / 0x5f89
     245 => std_logic_vector(to_unsigned(26738, 16)), -- 26738 / 0x6872
     246 => std_logic_vector(to_unsigned( 6030, 16)), --  6030 / 0x178e
     247 => std_logic_vector(to_unsigned(  505, 16)), --   505 / 0x01f9 -- last item of row
     248 => std_logic_vector(to_unsigned(   85, 16)), --    85 / 0x0055
     249 => std_logic_vector(to_unsigned(30326, 16)), -- 30326 / 0x7676
     250 => std_logic_vector(to_unsigned(22298, 16)), -- 22298 / 0x571a
     251 => std_logic_vector(to_unsigned(27562, 16)), -- 27562 / 0x6baa
     252 => std_logic_vector(to_unsigned(20131, 16)), -- 20131 / 0x4ea3
     253 => std_logic_vector(to_unsigned(26390, 16)), -- 26390 / 0x6716
     254 => std_logic_vector(to_unsigned( 6247, 16)), --  6247 / 0x1867
     255 => std_logic_vector(to_unsigned(24791, 16)), -- 24791 / 0x60d7 -- last item of row
     256 => std_logic_vector(to_unsigned(   86, 16)), --    86 / 0x0056
     257 => std_logic_vector(to_unsigned(  928, 16)), --   928 / 0x03a0
     258 => std_logic_vector(to_unsigned(29246, 16)), -- 29246 / 0x723e
     259 => std_logic_vector(to_unsigned(21246, 16)), -- 21246 / 0x52fe
     260 => std_logic_vector(to_unsigned(12400, 16)), -- 12400 / 0x3070
     261 => std_logic_vector(to_unsigned(15311, 16)), -- 15311 / 0x3bcf
     262 => std_logic_vector(to_unsigned(32309, 16)), -- 32309 / 0x7e35
     263 => std_logic_vector(to_unsigned(18608, 16)), -- 18608 / 0x48b0 -- last item of row
     264 => std_logic_vector(to_unsigned(   87, 16)), --    87 / 0x0057
     265 => std_logic_vector(to_unsigned(20314, 16)), -- 20314 / 0x4f5a
     266 => std_logic_vector(to_unsigned( 6025, 16)), --  6025 / 0x1789
     267 => std_logic_vector(to_unsigned(26689, 16)), -- 26689 / 0x6841
     268 => std_logic_vector(to_unsigned(16302, 16)), -- 16302 / 0x3fae
     269 => std_logic_vector(to_unsigned( 2296, 16)), --  2296 / 0x08f8
     270 => std_logic_vector(to_unsigned( 3244, 16)), --  3244 / 0x0cac
     271 => std_logic_vector(to_unsigned(19613, 16)), -- 19613 / 0x4c9d -- last item of row
     272 => std_logic_vector(to_unsigned(   88, 16)), --    88 / 0x0058
     273 => std_logic_vector(to_unsigned( 6237, 16)), --  6237 / 0x185d
     274 => std_logic_vector(to_unsigned(11943, 16)), -- 11943 / 0x2ea7
     275 => std_logic_vector(to_unsigned(22851, 16)), -- 22851 / 0x5943
     276 => std_logic_vector(to_unsigned(15642, 16)), -- 15642 / 0x3d1a
     277 => std_logic_vector(to_unsigned(23857, 16)), -- 23857 / 0x5d31
     278 => std_logic_vector(to_unsigned(15112, 16)), -- 15112 / 0x3b08
     279 => std_logic_vector(to_unsigned(20947, 16)), -- 20947 / 0x51d3 -- last item of row
     280 => std_logic_vector(to_unsigned(   89, 16)), --    89 / 0x0059
     281 => std_logic_vector(to_unsigned(26403, 16)), -- 26403 / 0x6723
     282 => std_logic_vector(to_unsigned(25168, 16)), -- 25168 / 0x6250
     283 => std_logic_vector(to_unsigned(19038, 16)), -- 19038 / 0x4a5e
     284 => std_logic_vector(to_unsigned(18384, 16)), -- 18384 / 0x47d0
     285 => std_logic_vector(to_unsigned( 8882, 16)), --  8882 / 0x22b2
     286 => std_logic_vector(to_unsigned(12719, 16)), -- 12719 / 0x31af
     287 => std_logic_vector(to_unsigned( 7093, 16)), --  7093 / 0x1bb5 -- last item of row
     288 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
     289 => std_logic_vector(to_unsigned(14567, 16)), -- 14567 / 0x38e7
     290 => std_logic_vector(to_unsigned(24965, 16)), -- 24965 / 0x6185 -- last item of row
     291 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
     292 => std_logic_vector(to_unsigned( 3908, 16)), --  3908 / 0x0f44
     293 => std_logic_vector(to_unsigned(  100, 16)), --   100 / 0x0064 -- last item of row
     294 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
     295 => std_logic_vector(to_unsigned(10279, 16)), -- 10279 / 0x2827
     296 => std_logic_vector(to_unsigned(  240, 16)), --   240 / 0x00f0 -- last item of row
     297 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
     298 => std_logic_vector(to_unsigned(24102, 16)), -- 24102 / 0x5e26
     299 => std_logic_vector(to_unsigned(  764, 16)), --   764 / 0x02fc -- last item of row
     300 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
     301 => std_logic_vector(to_unsigned(12383, 16)), -- 12383 / 0x305f
     302 => std_logic_vector(to_unsigned( 4173, 16)), --  4173 / 0x104d -- last item of row
     303 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
     304 => std_logic_vector(to_unsigned(13861, 16)), -- 13861 / 0x3625
     305 => std_logic_vector(to_unsigned(15918, 16)), -- 15918 / 0x3e2e -- last item of row
     306 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
     307 => std_logic_vector(to_unsigned(21327, 16)), -- 21327 / 0x534f
     308 => std_logic_vector(to_unsigned( 1046, 16)), --  1046 / 0x0416 -- last item of row
     309 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
     310 => std_logic_vector(to_unsigned( 5288, 16)), --  5288 / 0x14a8
     311 => std_logic_vector(to_unsigned(14579, 16)), -- 14579 / 0x38f3 -- last item of row
     312 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
     313 => std_logic_vector(to_unsigned(28158, 16)), -- 28158 / 0x6dfe
     314 => std_logic_vector(to_unsigned( 8069, 16)), --  8069 / 0x1f85 -- last item of row
     315 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
     316 => std_logic_vector(to_unsigned(16583, 16)), -- 16583 / 0x40c7
     317 => std_logic_vector(to_unsigned(11098, 16)), -- 11098 / 0x2b5a -- last item of row
     318 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
     319 => std_logic_vector(to_unsigned(16681, 16)), -- 16681 / 0x4129
     320 => std_logic_vector(to_unsigned(28363, 16)), -- 28363 / 0x6ecb -- last item of row
     321 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
     322 => std_logic_vector(to_unsigned(13980, 16)), -- 13980 / 0x369c
     323 => std_logic_vector(to_unsigned(24725, 16)), -- 24725 / 0x6095 -- last item of row
     324 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
     325 => std_logic_vector(to_unsigned(32169, 16)), -- 32169 / 0x7da9
     326 => std_logic_vector(to_unsigned(17989, 16)), -- 17989 / 0x4645 -- last item of row
     327 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
     328 => std_logic_vector(to_unsigned(10907, 16)), -- 10907 / 0x2a9b
     329 => std_logic_vector(to_unsigned( 2767, 16)), --  2767 / 0x0acf -- last item of row
     330 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
     331 => std_logic_vector(to_unsigned(21557, 16)), -- 21557 / 0x5435
     332 => std_logic_vector(to_unsigned( 3818, 16)), --  3818 / 0x0eea -- last item of row
     333 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
     334 => std_logic_vector(to_unsigned(26676, 16)), -- 26676 / 0x6834
     335 => std_logic_vector(to_unsigned(12422, 16)), -- 12422 / 0x3086 -- last item of row
     336 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
     337 => std_logic_vector(to_unsigned( 7676, 16)), --  7676 / 0x1dfc
     338 => std_logic_vector(to_unsigned( 8754, 16)), --  8754 / 0x2232 -- last item of row
     339 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
     340 => std_logic_vector(to_unsigned(14905, 16)), -- 14905 / 0x3a39
     341 => std_logic_vector(to_unsigned(20232, 16)), -- 20232 / 0x4f08 -- last item of row
     342 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
     343 => std_logic_vector(to_unsigned(15719, 16)), -- 15719 / 0x3d67
     344 => std_logic_vector(to_unsigned(24646, 16)), -- 24646 / 0x6046 -- last item of row
     345 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
     346 => std_logic_vector(to_unsigned(31942, 16)), -- 31942 / 0x7cc6
     347 => std_logic_vector(to_unsigned( 8589, 16)), --  8589 / 0x218d -- last item of row
     348 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
     349 => std_logic_vector(to_unsigned(19978, 16)), -- 19978 / 0x4e0a
     350 => std_logic_vector(to_unsigned(27197, 16)), -- 27197 / 0x6a3d -- last item of row
     351 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
     352 => std_logic_vector(to_unsigned(27060, 16)), -- 27060 / 0x69b4
     353 => std_logic_vector(to_unsigned(15071, 16)), -- 15071 / 0x3adf -- last item of row
     354 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
     355 => std_logic_vector(to_unsigned( 6071, 16)), --  6071 / 0x17b7
     356 => std_logic_vector(to_unsigned(26649, 16)), -- 26649 / 0x6819 -- last item of row
     357 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
     358 => std_logic_vector(to_unsigned(10393, 16)), -- 10393 / 0x2899
     359 => std_logic_vector(to_unsigned(11176, 16)), -- 11176 / 0x2ba8 -- last item of row
     360 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
     361 => std_logic_vector(to_unsigned( 9597, 16)), --  9597 / 0x257d
     362 => std_logic_vector(to_unsigned(13370, 16)), -- 13370 / 0x343a -- last item of row
     363 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
     364 => std_logic_vector(to_unsigned( 7081, 16)), --  7081 / 0x1ba9
     365 => std_logic_vector(to_unsigned(17677, 16)), -- 17677 / 0x450d -- last item of row
     366 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
     367 => std_logic_vector(to_unsigned( 1433, 16)), --  1433 / 0x0599
     368 => std_logic_vector(to_unsigned(19513, 16)), -- 19513 / 0x4c39 -- last item of row
     369 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
     370 => std_logic_vector(to_unsigned(26925, 16)), -- 26925 / 0x692d
     371 => std_logic_vector(to_unsigned( 9014, 16)), --  9014 / 0x2336 -- last item of row
     372 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
     373 => std_logic_vector(to_unsigned(19202, 16)), -- 19202 / 0x4b02
     374 => std_logic_vector(to_unsigned( 8900, 16)), --  8900 / 0x22c4 -- last item of row
     375 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
     376 => std_logic_vector(to_unsigned(18152, 16)), -- 18152 / 0x46e8
     377 => std_logic_vector(to_unsigned(30647, 16)), -- 30647 / 0x77b7 -- last item of row
     378 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
     379 => std_logic_vector(to_unsigned(20803, 16)), -- 20803 / 0x5143
     380 => std_logic_vector(to_unsigned( 1737, 16)), --  1737 / 0x06c9 -- last item of row
     381 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
     382 => std_logic_vector(to_unsigned(11804, 16)), -- 11804 / 0x2e1c
     383 => std_logic_vector(to_unsigned(25221, 16)), -- 25221 / 0x6285 -- last item of row
     384 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
     385 => std_logic_vector(to_unsigned(31683, 16)), -- 31683 / 0x7bc3
     386 => std_logic_vector(to_unsigned(17783, 16)), -- 17783 / 0x4577 -- last item of row
     387 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
     388 => std_logic_vector(to_unsigned(29694, 16)), -- 29694 / 0x73fe
     389 => std_logic_vector(to_unsigned( 9345, 16)), --  9345 / 0x2481 -- last item of row
     390 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
     391 => std_logic_vector(to_unsigned(12280, 16)), -- 12280 / 0x2ff8
     392 => std_logic_vector(to_unsigned(26611, 16)), -- 26611 / 0x67f3 -- last item of row
     393 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
     394 => std_logic_vector(to_unsigned( 6526, 16)), --  6526 / 0x197e
     395 => std_logic_vector(to_unsigned(26122, 16)), -- 26122 / 0x660a -- last item of row
     396 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
     397 => std_logic_vector(to_unsigned(26165, 16)), -- 26165 / 0x6635
     398 => std_logic_vector(to_unsigned(11241, 16)), -- 11241 / 0x2be9 -- last item of row
     399 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
     400 => std_logic_vector(to_unsigned( 7666, 16)), --  7666 / 0x1df2
     401 => std_logic_vector(to_unsigned(26962, 16)), -- 26962 / 0x6952 -- last item of row
     402 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
     403 => std_logic_vector(to_unsigned(16290, 16)), -- 16290 / 0x3fa2
     404 => std_logic_vector(to_unsigned( 8480, 16)), --  8480 / 0x2120 -- last item of row
     405 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
     406 => std_logic_vector(to_unsigned(11774, 16)), -- 11774 / 0x2dfe
     407 => std_logic_vector(to_unsigned(10120, 16)), -- 10120 / 0x2788 -- last item of row
     408 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
     409 => std_logic_vector(to_unsigned(30051, 16)), -- 30051 / 0x7563
     410 => std_logic_vector(to_unsigned(30426, 16)), -- 30426 / 0x76da -- last item of row
     411 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
     412 => std_logic_vector(to_unsigned( 1335, 16)), --  1335 / 0x0537
     413 => std_logic_vector(to_unsigned(15424, 16)), -- 15424 / 0x3c40 -- last item of row
     414 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
     415 => std_logic_vector(to_unsigned( 6865, 16)), --  6865 / 0x1ad1
     416 => std_logic_vector(to_unsigned(17742, 16)), -- 17742 / 0x454e -- last item of row
     417 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
     418 => std_logic_vector(to_unsigned(31779, 16)), -- 31779 / 0x7c23
     419 => std_logic_vector(to_unsigned(12489, 16)), -- 12489 / 0x30c9 -- last item of row
     420 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
     421 => std_logic_vector(to_unsigned(32120, 16)), -- 32120 / 0x7d78
     422 => std_logic_vector(to_unsigned(21001, 16)), -- 21001 / 0x5209 -- last item of row
     423 => std_logic_vector(to_unsigned(   45, 16)), --    45 / 0x002d
     424 => std_logic_vector(to_unsigned(14508, 16)), -- 14508 / 0x38ac
     425 => std_logic_vector(to_unsigned( 6996, 16)), --  6996 / 0x1b54 -- last item of row
     426 => std_logic_vector(to_unsigned(   46, 16)), --    46 / 0x002e
     427 => std_logic_vector(to_unsigned(  979, 16)), --   979 / 0x03d3
     428 => std_logic_vector(to_unsigned(25024, 16)), -- 25024 / 0x61c0 -- last item of row
     429 => std_logic_vector(to_unsigned(   47, 16)), --    47 / 0x002f
     430 => std_logic_vector(to_unsigned( 4554, 16)), --  4554 / 0x11ca
     431 => std_logic_vector(to_unsigned(21896, 16)), -- 21896 / 0x5588 -- last item of row
     432 => std_logic_vector(to_unsigned(   48, 16)), --    48 / 0x0030
     433 => std_logic_vector(to_unsigned( 7989, 16)), --  7989 / 0x1f35
     434 => std_logic_vector(to_unsigned(21777, 16)), -- 21777 / 0x5511 -- last item of row
     435 => std_logic_vector(to_unsigned(   49, 16)), --    49 / 0x0031
     436 => std_logic_vector(to_unsigned( 4972, 16)), --  4972 / 0x136c
     437 => std_logic_vector(to_unsigned(20661, 16)), -- 20661 / 0x50b5 -- last item of row
     438 => std_logic_vector(to_unsigned(   50, 16)), --    50 / 0x0032
     439 => std_logic_vector(to_unsigned( 6612, 16)), --  6612 / 0x19d4
     440 => std_logic_vector(to_unsigned( 2730, 16)), --  2730 / 0x0aaa -- last item of row
     441 => std_logic_vector(to_unsigned(   51, 16)), --    51 / 0x0033
     442 => std_logic_vector(to_unsigned(12742, 16)), -- 12742 / 0x31c6
     443 => std_logic_vector(to_unsigned( 4418, 16)), --  4418 / 0x1142 -- last item of row
     444 => std_logic_vector(to_unsigned(   52, 16)), --    52 / 0x0034
     445 => std_logic_vector(to_unsigned(29194, 16)), -- 29194 / 0x720a
     446 => std_logic_vector(to_unsigned(  595, 16)), --   595 / 0x0253 -- last item of row
     447 => std_logic_vector(to_unsigned(   53, 16)), --    53 / 0x0035
     448 => std_logic_vector(to_unsigned(19267, 16)), -- 19267 / 0x4b43
     449 => std_logic_vector(to_unsigned(20113, 16)), -- 20113 / 0x4e91 -- last item of row
    -- Table for fecframe_normal, C1_3
     450 => std_logic_vector(to_unsigned(34903, 16)), -- 34903 / 0x8857
     451 => std_logic_vector(to_unsigned(20927, 16)), -- 20927 / 0x51bf
     452 => std_logic_vector(to_unsigned(32093, 16)), -- 32093 / 0x7d5d
     453 => std_logic_vector(to_unsigned( 1052, 16)), --  1052 / 0x041c
     454 => std_logic_vector(to_unsigned(25611, 16)), -- 25611 / 0x640b
     455 => std_logic_vector(to_unsigned(16093, 16)), -- 16093 / 0x3edd
     456 => std_logic_vector(to_unsigned(16454, 16)), -- 16454 / 0x4046
     457 => std_logic_vector(to_unsigned( 5520, 16)), --  5520 / 0x1590
     458 => std_logic_vector(to_unsigned(  506, 16)), --   506 / 0x01fa
     459 => std_logic_vector(to_unsigned(37399, 16)), -- 37399 / 0x9217
     460 => std_logic_vector(to_unsigned(18518, 16)), -- 18518 / 0x4856
     461 => std_logic_vector(to_unsigned(21120, 16)), -- 21120 / 0x5280 -- last item of row
     462 => std_logic_vector(to_unsigned(11636, 16)), -- 11636 / 0x2d74
     463 => std_logic_vector(to_unsigned(14594, 16)), -- 14594 / 0x3902
     464 => std_logic_vector(to_unsigned(22158, 16)), -- 22158 / 0x568e
     465 => std_logic_vector(to_unsigned(14763, 16)), -- 14763 / 0x39ab
     466 => std_logic_vector(to_unsigned(15333, 16)), -- 15333 / 0x3be5
     467 => std_logic_vector(to_unsigned( 6838, 16)), --  6838 / 0x1ab6
     468 => std_logic_vector(to_unsigned(22222, 16)), -- 22222 / 0x56ce
     469 => std_logic_vector(to_unsigned(37856, 16)), -- 37856 / 0x93e0
     470 => std_logic_vector(to_unsigned(14985, 16)), -- 14985 / 0x3a89
     471 => std_logic_vector(to_unsigned(31041, 16)), -- 31041 / 0x7941
     472 => std_logic_vector(to_unsigned(18704, 16)), -- 18704 / 0x4910
     473 => std_logic_vector(to_unsigned(32910, 16)), -- 32910 / 0x808e -- last item of row
     474 => std_logic_vector(to_unsigned(17449, 16)), -- 17449 / 0x4429
     475 => std_logic_vector(to_unsigned( 1665, 16)), --  1665 / 0x0681
     476 => std_logic_vector(to_unsigned(35639, 16)), -- 35639 / 0x8b37
     477 => std_logic_vector(to_unsigned(16624, 16)), -- 16624 / 0x40f0
     478 => std_logic_vector(to_unsigned(12867, 16)), -- 12867 / 0x3243
     479 => std_logic_vector(to_unsigned(12449, 16)), -- 12449 / 0x30a1
     480 => std_logic_vector(to_unsigned(10241, 16)), -- 10241 / 0x2801
     481 => std_logic_vector(to_unsigned(11650, 16)), -- 11650 / 0x2d82
     482 => std_logic_vector(to_unsigned(25622, 16)), -- 25622 / 0x6416
     483 => std_logic_vector(to_unsigned(34372, 16)), -- 34372 / 0x8644
     484 => std_logic_vector(to_unsigned(19878, 16)), -- 19878 / 0x4da6
     485 => std_logic_vector(to_unsigned(26894, 16)), -- 26894 / 0x690e -- last item of row
     486 => std_logic_vector(to_unsigned(29235, 16)), -- 29235 / 0x7233
     487 => std_logic_vector(to_unsigned(19780, 16)), -- 19780 / 0x4d44
     488 => std_logic_vector(to_unsigned(36056, 16)), -- 36056 / 0x8cd8
     489 => std_logic_vector(to_unsigned(20129, 16)), -- 20129 / 0x4ea1
     490 => std_logic_vector(to_unsigned(20029, 16)), -- 20029 / 0x4e3d
     491 => std_logic_vector(to_unsigned( 5457, 16)), --  5457 / 0x1551
     492 => std_logic_vector(to_unsigned( 8157, 16)), --  8157 / 0x1fdd
     493 => std_logic_vector(to_unsigned(35554, 16)), -- 35554 / 0x8ae2
     494 => std_logic_vector(to_unsigned(21237, 16)), -- 21237 / 0x52f5
     495 => std_logic_vector(to_unsigned( 7943, 16)), --  7943 / 0x1f07
     496 => std_logic_vector(to_unsigned(13873, 16)), -- 13873 / 0x3631
     497 => std_logic_vector(to_unsigned(14980, 16)), -- 14980 / 0x3a84 -- last item of row
     498 => std_logic_vector(to_unsigned( 9912, 16)), --  9912 / 0x26b8
     499 => std_logic_vector(to_unsigned( 7143, 16)), --  7143 / 0x1be7
     500 => std_logic_vector(to_unsigned(35911, 16)), -- 35911 / 0x8c47
     501 => std_logic_vector(to_unsigned(12043, 16)), -- 12043 / 0x2f0b
     502 => std_logic_vector(to_unsigned(17360, 16)), -- 17360 / 0x43d0
     503 => std_logic_vector(to_unsigned(37253, 16)), -- 37253 / 0x9185
     504 => std_logic_vector(to_unsigned(25588, 16)), -- 25588 / 0x63f4
     505 => std_logic_vector(to_unsigned(11827, 16)), -- 11827 / 0x2e33
     506 => std_logic_vector(to_unsigned(29152, 16)), -- 29152 / 0x71e0
     507 => std_logic_vector(to_unsigned(21936, 16)), -- 21936 / 0x55b0
     508 => std_logic_vector(to_unsigned(24125, 16)), -- 24125 / 0x5e3d
     509 => std_logic_vector(to_unsigned(40870, 16)), -- 40870 / 0x9fa6 -- last item of row
     510 => std_logic_vector(to_unsigned(40701, 16)), -- 40701 / 0x9efd
     511 => std_logic_vector(to_unsigned(36035, 16)), -- 36035 / 0x8cc3
     512 => std_logic_vector(to_unsigned(39556, 16)), -- 39556 / 0x9a84
     513 => std_logic_vector(to_unsigned(12366, 16)), -- 12366 / 0x304e
     514 => std_logic_vector(to_unsigned(19946, 16)), -- 19946 / 0x4dea
     515 => std_logic_vector(to_unsigned(29072, 16)), -- 29072 / 0x7190
     516 => std_logic_vector(to_unsigned(16365, 16)), -- 16365 / 0x3fed
     517 => std_logic_vector(to_unsigned(35495, 16)), -- 35495 / 0x8aa7
     518 => std_logic_vector(to_unsigned(22686, 16)), -- 22686 / 0x589e
     519 => std_logic_vector(to_unsigned(11106, 16)), -- 11106 / 0x2b62
     520 => std_logic_vector(to_unsigned( 8756, 16)), --  8756 / 0x2234
     521 => std_logic_vector(to_unsigned(34863, 16)), -- 34863 / 0x882f -- last item of row
     522 => std_logic_vector(to_unsigned(19165, 16)), -- 19165 / 0x4add
     523 => std_logic_vector(to_unsigned(15702, 16)), -- 15702 / 0x3d56
     524 => std_logic_vector(to_unsigned(13536, 16)), -- 13536 / 0x34e0
     525 => std_logic_vector(to_unsigned(40238, 16)), -- 40238 / 0x9d2e
     526 => std_logic_vector(to_unsigned( 4465, 16)), --  4465 / 0x1171
     527 => std_logic_vector(to_unsigned(40034, 16)), -- 40034 / 0x9c62
     528 => std_logic_vector(to_unsigned(40590, 16)), -- 40590 / 0x9e8e
     529 => std_logic_vector(to_unsigned(37540, 16)), -- 37540 / 0x92a4
     530 => std_logic_vector(to_unsigned(17162, 16)), -- 17162 / 0x430a
     531 => std_logic_vector(to_unsigned( 1712, 16)), --  1712 / 0x06b0
     532 => std_logic_vector(to_unsigned(20577, 16)), -- 20577 / 0x5061
     533 => std_logic_vector(to_unsigned(14138, 16)), -- 14138 / 0x373a -- last item of row
     534 => std_logic_vector(to_unsigned(31338, 16)), -- 31338 / 0x7a6a
     535 => std_logic_vector(to_unsigned(19342, 16)), -- 19342 / 0x4b8e
     536 => std_logic_vector(to_unsigned( 9301, 16)), --  9301 / 0x2455
     537 => std_logic_vector(to_unsigned(39375, 16)), -- 39375 / 0x99cf
     538 => std_logic_vector(to_unsigned( 3211, 16)), --  3211 / 0x0c8b
     539 => std_logic_vector(to_unsigned( 1316, 16)), --  1316 / 0x0524
     540 => std_logic_vector(to_unsigned(33409, 16)), -- 33409 / 0x8281
     541 => std_logic_vector(to_unsigned(28670, 16)), -- 28670 / 0x6ffe
     542 => std_logic_vector(to_unsigned(12282, 16)), -- 12282 / 0x2ffa
     543 => std_logic_vector(to_unsigned( 6118, 16)), --  6118 / 0x17e6
     544 => std_logic_vector(to_unsigned(29236, 16)), -- 29236 / 0x7234
     545 => std_logic_vector(to_unsigned(35787, 16)), -- 35787 / 0x8bcb -- last item of row
     546 => std_logic_vector(to_unsigned(11504, 16)), -- 11504 / 0x2cf0
     547 => std_logic_vector(to_unsigned(30506, 16)), -- 30506 / 0x772a
     548 => std_logic_vector(to_unsigned(19558, 16)), -- 19558 / 0x4c66
     549 => std_logic_vector(to_unsigned( 5100, 16)), --  5100 / 0x13ec
     550 => std_logic_vector(to_unsigned(24188, 16)), -- 24188 / 0x5e7c
     551 => std_logic_vector(to_unsigned(24738, 16)), -- 24738 / 0x60a2
     552 => std_logic_vector(to_unsigned(30397, 16)), -- 30397 / 0x76bd
     553 => std_logic_vector(to_unsigned(33775, 16)), -- 33775 / 0x83ef
     554 => std_logic_vector(to_unsigned( 9699, 16)), --  9699 / 0x25e3
     555 => std_logic_vector(to_unsigned( 6215, 16)), --  6215 / 0x1847
     556 => std_logic_vector(to_unsigned( 3397, 16)), --  3397 / 0x0d45
     557 => std_logic_vector(to_unsigned(37451, 16)), -- 37451 / 0x924b -- last item of row
     558 => std_logic_vector(to_unsigned(34689, 16)), -- 34689 / 0x8781
     559 => std_logic_vector(to_unsigned(23126, 16)), -- 23126 / 0x5a56
     560 => std_logic_vector(to_unsigned( 7571, 16)), --  7571 / 0x1d93
     561 => std_logic_vector(to_unsigned( 1058, 16)), --  1058 / 0x0422
     562 => std_logic_vector(to_unsigned(12127, 16)), -- 12127 / 0x2f5f
     563 => std_logic_vector(to_unsigned(27518, 16)), -- 27518 / 0x6b7e
     564 => std_logic_vector(to_unsigned(23064, 16)), -- 23064 / 0x5a18
     565 => std_logic_vector(to_unsigned(11265, 16)), -- 11265 / 0x2c01
     566 => std_logic_vector(to_unsigned(14867, 16)), -- 14867 / 0x3a13
     567 => std_logic_vector(to_unsigned(30451, 16)), -- 30451 / 0x76f3
     568 => std_logic_vector(to_unsigned(28289, 16)), -- 28289 / 0x6e81
     569 => std_logic_vector(to_unsigned( 2966, 16)), --  2966 / 0x0b96 -- last item of row
     570 => std_logic_vector(to_unsigned(11660, 16)), -- 11660 / 0x2d8c
     571 => std_logic_vector(to_unsigned(15334, 16)), -- 15334 / 0x3be6
     572 => std_logic_vector(to_unsigned(16867, 16)), -- 16867 / 0x41e3
     573 => std_logic_vector(to_unsigned(15160, 16)), -- 15160 / 0x3b38
     574 => std_logic_vector(to_unsigned(38343, 16)), -- 38343 / 0x95c7
     575 => std_logic_vector(to_unsigned( 3778, 16)), --  3778 / 0x0ec2
     576 => std_logic_vector(to_unsigned( 4265, 16)), --  4265 / 0x10a9
     577 => std_logic_vector(to_unsigned(39139, 16)), -- 39139 / 0x98e3
     578 => std_logic_vector(to_unsigned(17293, 16)), -- 17293 / 0x438d
     579 => std_logic_vector(to_unsigned(26229, 16)), -- 26229 / 0x6675
     580 => std_logic_vector(to_unsigned(42604, 16)), -- 42604 / 0xa66c
     581 => std_logic_vector(to_unsigned(13486, 16)), -- 13486 / 0x34ae -- last item of row
     582 => std_logic_vector(to_unsigned(31497, 16)), -- 31497 / 0x7b09
     583 => std_logic_vector(to_unsigned( 1365, 16)), --  1365 / 0x0555
     584 => std_logic_vector(to_unsigned(14828, 16)), -- 14828 / 0x39ec
     585 => std_logic_vector(to_unsigned( 7453, 16)), --  7453 / 0x1d1d
     586 => std_logic_vector(to_unsigned(26350, 16)), -- 26350 / 0x66ee
     587 => std_logic_vector(to_unsigned(41346, 16)), -- 41346 / 0xa182
     588 => std_logic_vector(to_unsigned(28643, 16)), -- 28643 / 0x6fe3
     589 => std_logic_vector(to_unsigned(23421, 16)), -- 23421 / 0x5b7d
     590 => std_logic_vector(to_unsigned( 8354, 16)), --  8354 / 0x20a2
     591 => std_logic_vector(to_unsigned(16255, 16)), -- 16255 / 0x3f7f
     592 => std_logic_vector(to_unsigned(11055, 16)), -- 11055 / 0x2b2f
     593 => std_logic_vector(to_unsigned(24279, 16)), -- 24279 / 0x5ed7 -- last item of row
     594 => std_logic_vector(to_unsigned(15687, 16)), -- 15687 / 0x3d47
     595 => std_logic_vector(to_unsigned(12467, 16)), -- 12467 / 0x30b3
     596 => std_logic_vector(to_unsigned(13906, 16)), -- 13906 / 0x3652
     597 => std_logic_vector(to_unsigned( 5215, 16)), --  5215 / 0x145f
     598 => std_logic_vector(to_unsigned(41328, 16)), -- 41328 / 0xa170
     599 => std_logic_vector(to_unsigned(23755, 16)), -- 23755 / 0x5ccb
     600 => std_logic_vector(to_unsigned(20800, 16)), -- 20800 / 0x5140
     601 => std_logic_vector(to_unsigned( 6447, 16)), --  6447 / 0x192f
     602 => std_logic_vector(to_unsigned( 7970, 16)), --  7970 / 0x1f22
     603 => std_logic_vector(to_unsigned( 2803, 16)), --  2803 / 0x0af3
     604 => std_logic_vector(to_unsigned(33262, 16)), -- 33262 / 0x81ee
     605 => std_logic_vector(to_unsigned(39843, 16)), -- 39843 / 0x9ba3 -- last item of row
     606 => std_logic_vector(to_unsigned( 5363, 16)), --  5363 / 0x14f3
     607 => std_logic_vector(to_unsigned(22469, 16)), -- 22469 / 0x57c5
     608 => std_logic_vector(to_unsigned(38091, 16)), -- 38091 / 0x94cb
     609 => std_logic_vector(to_unsigned(28457, 16)), -- 28457 / 0x6f29
     610 => std_logic_vector(to_unsigned(36696, 16)), -- 36696 / 0x8f58
     611 => std_logic_vector(to_unsigned(34471, 16)), -- 34471 / 0x86a7
     612 => std_logic_vector(to_unsigned(23619, 16)), -- 23619 / 0x5c43
     613 => std_logic_vector(to_unsigned( 2404, 16)), --  2404 / 0x0964
     614 => std_logic_vector(to_unsigned(24229, 16)), -- 24229 / 0x5ea5
     615 => std_logic_vector(to_unsigned(41754, 16)), -- 41754 / 0xa31a
     616 => std_logic_vector(to_unsigned( 1297, 16)), --  1297 / 0x0511
     617 => std_logic_vector(to_unsigned(18563, 16)), -- 18563 / 0x4883 -- last item of row
     618 => std_logic_vector(to_unsigned( 3673, 16)), --  3673 / 0x0e59
     619 => std_logic_vector(to_unsigned(39070, 16)), -- 39070 / 0x989e
     620 => std_logic_vector(to_unsigned(14480, 16)), -- 14480 / 0x3890
     621 => std_logic_vector(to_unsigned(30279, 16)), -- 30279 / 0x7647
     622 => std_logic_vector(to_unsigned(37483, 16)), -- 37483 / 0x926b
     623 => std_logic_vector(to_unsigned( 7580, 16)), --  7580 / 0x1d9c
     624 => std_logic_vector(to_unsigned(29519, 16)), -- 29519 / 0x734f
     625 => std_logic_vector(to_unsigned(30519, 16)), -- 30519 / 0x7737
     626 => std_logic_vector(to_unsigned(39831, 16)), -- 39831 / 0x9b97
     627 => std_logic_vector(to_unsigned(20252, 16)), -- 20252 / 0x4f1c
     628 => std_logic_vector(to_unsigned(18132, 16)), -- 18132 / 0x46d4
     629 => std_logic_vector(to_unsigned(20010, 16)), -- 20010 / 0x4e2a -- last item of row
     630 => std_logic_vector(to_unsigned(34386, 16)), -- 34386 / 0x8652
     631 => std_logic_vector(to_unsigned( 7252, 16)), --  7252 / 0x1c54
     632 => std_logic_vector(to_unsigned(27526, 16)), -- 27526 / 0x6b86
     633 => std_logic_vector(to_unsigned(12950, 16)), -- 12950 / 0x3296
     634 => std_logic_vector(to_unsigned( 6875, 16)), --  6875 / 0x1adb
     635 => std_logic_vector(to_unsigned(43020, 16)), -- 43020 / 0xa80c
     636 => std_logic_vector(to_unsigned(31566, 16)), -- 31566 / 0x7b4e
     637 => std_logic_vector(to_unsigned(39069, 16)), -- 39069 / 0x989d
     638 => std_logic_vector(to_unsigned(18985, 16)), -- 18985 / 0x4a29
     639 => std_logic_vector(to_unsigned(15541, 16)), -- 15541 / 0x3cb5
     640 => std_logic_vector(to_unsigned(40020, 16)), -- 40020 / 0x9c54
     641 => std_logic_vector(to_unsigned(16715, 16)), -- 16715 / 0x414b -- last item of row
     642 => std_logic_vector(to_unsigned( 1721, 16)), --  1721 / 0x06b9
     643 => std_logic_vector(to_unsigned(37332, 16)), -- 37332 / 0x91d4
     644 => std_logic_vector(to_unsigned(39953, 16)), -- 39953 / 0x9c11
     645 => std_logic_vector(to_unsigned(17430, 16)), -- 17430 / 0x4416
     646 => std_logic_vector(to_unsigned(32134, 16)), -- 32134 / 0x7d86
     647 => std_logic_vector(to_unsigned(29162, 16)), -- 29162 / 0x71ea
     648 => std_logic_vector(to_unsigned(10490, 16)), -- 10490 / 0x28fa
     649 => std_logic_vector(to_unsigned(12971, 16)), -- 12971 / 0x32ab
     650 => std_logic_vector(to_unsigned(28581, 16)), -- 28581 / 0x6fa5
     651 => std_logic_vector(to_unsigned(29331, 16)), -- 29331 / 0x7293
     652 => std_logic_vector(to_unsigned( 6489, 16)), --  6489 / 0x1959
     653 => std_logic_vector(to_unsigned(35383, 16)), -- 35383 / 0x8a37 -- last item of row
     654 => std_logic_vector(to_unsigned(  736, 16)), --   736 / 0x02e0
     655 => std_logic_vector(to_unsigned( 7022, 16)), --  7022 / 0x1b6e
     656 => std_logic_vector(to_unsigned(42349, 16)), -- 42349 / 0xa56d
     657 => std_logic_vector(to_unsigned( 8783, 16)), --  8783 / 0x224f
     658 => std_logic_vector(to_unsigned( 6767, 16)), --  6767 / 0x1a6f
     659 => std_logic_vector(to_unsigned(11871, 16)), -- 11871 / 0x2e5f
     660 => std_logic_vector(to_unsigned(21675, 16)), -- 21675 / 0x54ab
     661 => std_logic_vector(to_unsigned(10325, 16)), -- 10325 / 0x2855
     662 => std_logic_vector(to_unsigned(11548, 16)), -- 11548 / 0x2d1c
     663 => std_logic_vector(to_unsigned(25978, 16)), -- 25978 / 0x657a
     664 => std_logic_vector(to_unsigned(  431, 16)), --   431 / 0x01af
     665 => std_logic_vector(to_unsigned(24085, 16)), -- 24085 / 0x5e15 -- last item of row
     666 => std_logic_vector(to_unsigned( 1925, 16)), --  1925 / 0x0785
     667 => std_logic_vector(to_unsigned(10602, 16)), -- 10602 / 0x296a
     668 => std_logic_vector(to_unsigned(28585, 16)), -- 28585 / 0x6fa9
     669 => std_logic_vector(to_unsigned(12170, 16)), -- 12170 / 0x2f8a
     670 => std_logic_vector(to_unsigned(15156, 16)), -- 15156 / 0x3b34
     671 => std_logic_vector(to_unsigned(34404, 16)), -- 34404 / 0x8664
     672 => std_logic_vector(to_unsigned( 8351, 16)), --  8351 / 0x209f
     673 => std_logic_vector(to_unsigned(13273, 16)), -- 13273 / 0x33d9
     674 => std_logic_vector(to_unsigned(20208, 16)), -- 20208 / 0x4ef0
     675 => std_logic_vector(to_unsigned( 5800, 16)), --  5800 / 0x16a8
     676 => std_logic_vector(to_unsigned(15367, 16)), -- 15367 / 0x3c07
     677 => std_logic_vector(to_unsigned(21764, 16)), -- 21764 / 0x5504 -- last item of row
     678 => std_logic_vector(to_unsigned(16279, 16)), -- 16279 / 0x3f97
     679 => std_logic_vector(to_unsigned(37832, 16)), -- 37832 / 0x93c8
     680 => std_logic_vector(to_unsigned(34792, 16)), -- 34792 / 0x87e8
     681 => std_logic_vector(to_unsigned(21250, 16)), -- 21250 / 0x5302
     682 => std_logic_vector(to_unsigned(34192, 16)), -- 34192 / 0x8590
     683 => std_logic_vector(to_unsigned( 7406, 16)), --  7406 / 0x1cee
     684 => std_logic_vector(to_unsigned(41488, 16)), -- 41488 / 0xa210
     685 => std_logic_vector(to_unsigned(18346, 16)), -- 18346 / 0x47aa
     686 => std_logic_vector(to_unsigned(29227, 16)), -- 29227 / 0x722b
     687 => std_logic_vector(to_unsigned(26127, 16)), -- 26127 / 0x660f
     688 => std_logic_vector(to_unsigned(25493, 16)), -- 25493 / 0x6395
     689 => std_logic_vector(to_unsigned( 7048, 16)), --  7048 / 0x1b88 -- last item of row
     690 => std_logic_vector(to_unsigned(39948, 16)), -- 39948 / 0x9c0c
     691 => std_logic_vector(to_unsigned(28229, 16)), -- 28229 / 0x6e45
     692 => std_logic_vector(to_unsigned(24899, 16)), -- 24899 / 0x6143 -- last item of row
     693 => std_logic_vector(to_unsigned(17408, 16)), -- 17408 / 0x4400
     694 => std_logic_vector(to_unsigned(14274, 16)), -- 14274 / 0x37c2
     695 => std_logic_vector(to_unsigned(38993, 16)), -- 38993 / 0x9851 -- last item of row
     696 => std_logic_vector(to_unsigned(38774, 16)), -- 38774 / 0x9776
     697 => std_logic_vector(to_unsigned(15968, 16)), -- 15968 / 0x3e60
     698 => std_logic_vector(to_unsigned(28459, 16)), -- 28459 / 0x6f2b -- last item of row
     699 => std_logic_vector(to_unsigned(41404, 16)), -- 41404 / 0xa1bc
     700 => std_logic_vector(to_unsigned(27249, 16)), -- 27249 / 0x6a71
     701 => std_logic_vector(to_unsigned(27425, 16)), -- 27425 / 0x6b21 -- last item of row
     702 => std_logic_vector(to_unsigned(41229, 16)), -- 41229 / 0xa10d
     703 => std_logic_vector(to_unsigned( 6082, 16)), --  6082 / 0x17c2
     704 => std_logic_vector(to_unsigned(43114, 16)), -- 43114 / 0xa86a -- last item of row
     705 => std_logic_vector(to_unsigned(13957, 16)), -- 13957 / 0x3685
     706 => std_logic_vector(to_unsigned( 4979, 16)), --  4979 / 0x1373
     707 => std_logic_vector(to_unsigned(40654, 16)), -- 40654 / 0x9ece -- last item of row
     708 => std_logic_vector(to_unsigned( 3093, 16)), --  3093 / 0x0c15
     709 => std_logic_vector(to_unsigned( 3438, 16)), --  3438 / 0x0d6e
     710 => std_logic_vector(to_unsigned(34992, 16)), -- 34992 / 0x88b0 -- last item of row
     711 => std_logic_vector(to_unsigned(34082, 16)), -- 34082 / 0x8522
     712 => std_logic_vector(to_unsigned( 6172, 16)), --  6172 / 0x181c
     713 => std_logic_vector(to_unsigned(28760, 16)), -- 28760 / 0x7058 -- last item of row
     714 => std_logic_vector(to_unsigned(42210, 16)), -- 42210 / 0xa4e2
     715 => std_logic_vector(to_unsigned(34141, 16)), -- 34141 / 0x855d
     716 => std_logic_vector(to_unsigned(41021, 16)), -- 41021 / 0xa03d -- last item of row
     717 => std_logic_vector(to_unsigned(14705, 16)), -- 14705 / 0x3971
     718 => std_logic_vector(to_unsigned(17783, 16)), -- 17783 / 0x4577
     719 => std_logic_vector(to_unsigned(10134, 16)), -- 10134 / 0x2796 -- last item of row
     720 => std_logic_vector(to_unsigned(41755, 16)), -- 41755 / 0xa31b
     721 => std_logic_vector(to_unsigned(39884, 16)), -- 39884 / 0x9bcc
     722 => std_logic_vector(to_unsigned(22773, 16)), -- 22773 / 0x58f5 -- last item of row
     723 => std_logic_vector(to_unsigned(14615, 16)), -- 14615 / 0x3917
     724 => std_logic_vector(to_unsigned(15593, 16)), -- 15593 / 0x3ce9
     725 => std_logic_vector(to_unsigned( 1642, 16)), --  1642 / 0x066a -- last item of row
     726 => std_logic_vector(to_unsigned(29111, 16)), -- 29111 / 0x71b7
     727 => std_logic_vector(to_unsigned(37061, 16)), -- 37061 / 0x90c5
     728 => std_logic_vector(to_unsigned(39860, 16)), -- 39860 / 0x9bb4 -- last item of row
     729 => std_logic_vector(to_unsigned( 9579, 16)), --  9579 / 0x256b
     730 => std_logic_vector(to_unsigned(33552, 16)), -- 33552 / 0x8310
     731 => std_logic_vector(to_unsigned(  633, 16)), --   633 / 0x0279 -- last item of row
     732 => std_logic_vector(to_unsigned(12951, 16)), -- 12951 / 0x3297
     733 => std_logic_vector(to_unsigned(21137, 16)), -- 21137 / 0x5291
     734 => std_logic_vector(to_unsigned(39608, 16)), -- 39608 / 0x9ab8 -- last item of row
     735 => std_logic_vector(to_unsigned(38244, 16)), -- 38244 / 0x9564
     736 => std_logic_vector(to_unsigned(27361, 16)), -- 27361 / 0x6ae1
     737 => std_logic_vector(to_unsigned(29417, 16)), -- 29417 / 0x72e9 -- last item of row
     738 => std_logic_vector(to_unsigned( 2939, 16)), --  2939 / 0x0b7b
     739 => std_logic_vector(to_unsigned(10172, 16)), -- 10172 / 0x27bc
     740 => std_logic_vector(to_unsigned(36479, 16)), -- 36479 / 0x8e7f -- last item of row
     741 => std_logic_vector(to_unsigned(29094, 16)), -- 29094 / 0x71a6
     742 => std_logic_vector(to_unsigned( 5357, 16)), --  5357 / 0x14ed
     743 => std_logic_vector(to_unsigned(19224, 16)), -- 19224 / 0x4b18 -- last item of row
     744 => std_logic_vector(to_unsigned( 9562, 16)), --  9562 / 0x255a
     745 => std_logic_vector(to_unsigned(24436, 16)), -- 24436 / 0x5f74
     746 => std_logic_vector(to_unsigned(28637, 16)), -- 28637 / 0x6fdd -- last item of row
     747 => std_logic_vector(to_unsigned(40177, 16)), -- 40177 / 0x9cf1
     748 => std_logic_vector(to_unsigned( 2326, 16)), --  2326 / 0x0916
     749 => std_logic_vector(to_unsigned(13504, 16)), -- 13504 / 0x34c0 -- last item of row
     750 => std_logic_vector(to_unsigned( 6834, 16)), --  6834 / 0x1ab2
     751 => std_logic_vector(to_unsigned(21583, 16)), -- 21583 / 0x544f
     752 => std_logic_vector(to_unsigned(42516, 16)), -- 42516 / 0xa614 -- last item of row
     753 => std_logic_vector(to_unsigned(40651, 16)), -- 40651 / 0x9ecb
     754 => std_logic_vector(to_unsigned(42810, 16)), -- 42810 / 0xa73a
     755 => std_logic_vector(to_unsigned(25709, 16)), -- 25709 / 0x646d -- last item of row
     756 => std_logic_vector(to_unsigned(31557, 16)), -- 31557 / 0x7b45
     757 => std_logic_vector(to_unsigned(32138, 16)), -- 32138 / 0x7d8a
     758 => std_logic_vector(to_unsigned(38142, 16)), -- 38142 / 0x94fe -- last item of row
     759 => std_logic_vector(to_unsigned(18624, 16)), -- 18624 / 0x48c0
     760 => std_logic_vector(to_unsigned(41867, 16)), -- 41867 / 0xa38b
     761 => std_logic_vector(to_unsigned(39296, 16)), -- 39296 / 0x9980 -- last item of row
     762 => std_logic_vector(to_unsigned(37560, 16)), -- 37560 / 0x92b8
     763 => std_logic_vector(to_unsigned(14295, 16)), -- 14295 / 0x37d7
     764 => std_logic_vector(to_unsigned(16245, 16)), -- 16245 / 0x3f75 -- last item of row
     765 => std_logic_vector(to_unsigned( 6821, 16)), --  6821 / 0x1aa5
     766 => std_logic_vector(to_unsigned(21679, 16)), -- 21679 / 0x54af
     767 => std_logic_vector(to_unsigned(31570, 16)), -- 31570 / 0x7b52 -- last item of row
     768 => std_logic_vector(to_unsigned(25339, 16)), -- 25339 / 0x62fb
     769 => std_logic_vector(to_unsigned(25083, 16)), -- 25083 / 0x61fb
     770 => std_logic_vector(to_unsigned(22081, 16)), -- 22081 / 0x5641 -- last item of row
     771 => std_logic_vector(to_unsigned( 8047, 16)), --  8047 / 0x1f6f
     772 => std_logic_vector(to_unsigned(  697, 16)), --   697 / 0x02b9
     773 => std_logic_vector(to_unsigned(35268, 16)), -- 35268 / 0x89c4 -- last item of row
     774 => std_logic_vector(to_unsigned( 9884, 16)), --  9884 / 0x269c
     775 => std_logic_vector(to_unsigned(17073, 16)), -- 17073 / 0x42b1
     776 => std_logic_vector(to_unsigned(19995, 16)), -- 19995 / 0x4e1b -- last item of row
     777 => std_logic_vector(to_unsigned(26848, 16)), -- 26848 / 0x68e0
     778 => std_logic_vector(to_unsigned(35245, 16)), -- 35245 / 0x89ad
     779 => std_logic_vector(to_unsigned( 8390, 16)), --  8390 / 0x20c6 -- last item of row
     780 => std_logic_vector(to_unsigned(18658, 16)), -- 18658 / 0x48e2
     781 => std_logic_vector(to_unsigned(16134, 16)), -- 16134 / 0x3f06
     782 => std_logic_vector(to_unsigned(14807, 16)), -- 14807 / 0x39d7 -- last item of row
     783 => std_logic_vector(to_unsigned(12201, 16)), -- 12201 / 0x2fa9
     784 => std_logic_vector(to_unsigned(32944, 16)), -- 32944 / 0x80b0
     785 => std_logic_vector(to_unsigned( 5035, 16)), --  5035 / 0x13ab -- last item of row
     786 => std_logic_vector(to_unsigned(25236, 16)), -- 25236 / 0x6294
     787 => std_logic_vector(to_unsigned( 1216, 16)), --  1216 / 0x04c0
     788 => std_logic_vector(to_unsigned(38986, 16)), -- 38986 / 0x984a -- last item of row
     789 => std_logic_vector(to_unsigned(42994, 16)), -- 42994 / 0xa7f2
     790 => std_logic_vector(to_unsigned(24782, 16)), -- 24782 / 0x60ce
     791 => std_logic_vector(to_unsigned( 8681, 16)), --  8681 / 0x21e9 -- last item of row
     792 => std_logic_vector(to_unsigned(28321, 16)), -- 28321 / 0x6ea1
     793 => std_logic_vector(to_unsigned( 4932, 16)), --  4932 / 0x1344
     794 => std_logic_vector(to_unsigned(34249, 16)), -- 34249 / 0x85c9 -- last item of row
     795 => std_logic_vector(to_unsigned( 4107, 16)), --  4107 / 0x100b
     796 => std_logic_vector(to_unsigned(29382, 16)), -- 29382 / 0x72c6
     797 => std_logic_vector(to_unsigned(32124, 16)), -- 32124 / 0x7d7c -- last item of row
     798 => std_logic_vector(to_unsigned(22157, 16)), -- 22157 / 0x568d
     799 => std_logic_vector(to_unsigned( 2624, 16)), --  2624 / 0x0a40
     800 => std_logic_vector(to_unsigned(14468, 16)), -- 14468 / 0x3884 -- last item of row
     801 => std_logic_vector(to_unsigned(38788, 16)), -- 38788 / 0x9784
     802 => std_logic_vector(to_unsigned(27081, 16)), -- 27081 / 0x69c9
     803 => std_logic_vector(to_unsigned( 7936, 16)), --  7936 / 0x1f00 -- last item of row
     804 => std_logic_vector(to_unsigned( 4368, 16)), --  4368 / 0x1110
     805 => std_logic_vector(to_unsigned(26148, 16)), -- 26148 / 0x6624
     806 => std_logic_vector(to_unsigned(10578, 16)), -- 10578 / 0x2952 -- last item of row
     807 => std_logic_vector(to_unsigned(25353, 16)), -- 25353 / 0x6309
     808 => std_logic_vector(to_unsigned( 4122, 16)), --  4122 / 0x101a
     809 => std_logic_vector(to_unsigned(39751, 16)), -- 39751 / 0x9b47 -- last item of row
    -- Table for fecframe_normal, C1_4
     810 => std_logic_vector(to_unsigned(23606, 16)), -- 23606 / 0x5c36
     811 => std_logic_vector(to_unsigned(36098, 16)), -- 36098 / 0x8d02
     812 => std_logic_vector(to_unsigned( 1140, 16)), --  1140 / 0x0474
     813 => std_logic_vector(to_unsigned(28859, 16)), -- 28859 / 0x70bb
     814 => std_logic_vector(to_unsigned(18148, 16)), -- 18148 / 0x46e4
     815 => std_logic_vector(to_unsigned(18510, 16)), -- 18510 / 0x484e
     816 => std_logic_vector(to_unsigned( 6226, 16)), --  6226 / 0x1852
     817 => std_logic_vector(to_unsigned(  540, 16)), --   540 / 0x021c
     818 => std_logic_vector(to_unsigned(42014, 16)), -- 42014 / 0xa41e
     819 => std_logic_vector(to_unsigned(20879, 16)), -- 20879 / 0x518f
     820 => std_logic_vector(to_unsigned(23802, 16)), -- 23802 / 0x5cfa
     821 => std_logic_vector(to_unsigned(47088, 16)), -- 47088 / 0xb7f0 -- last item of row
     822 => std_logic_vector(to_unsigned(16419, 16)), -- 16419 / 0x4023
     823 => std_logic_vector(to_unsigned(24928, 16)), -- 24928 / 0x6160
     824 => std_logic_vector(to_unsigned(16609, 16)), -- 16609 / 0x40e1
     825 => std_logic_vector(to_unsigned(17248, 16)), -- 17248 / 0x4360
     826 => std_logic_vector(to_unsigned( 7693, 16)), --  7693 / 0x1e0d
     827 => std_logic_vector(to_unsigned(24997, 16)), -- 24997 / 0x61a5
     828 => std_logic_vector(to_unsigned(42587, 16)), -- 42587 / 0xa65b
     829 => std_logic_vector(to_unsigned(16858, 16)), -- 16858 / 0x41da
     830 => std_logic_vector(to_unsigned(34921, 16)), -- 34921 / 0x8869
     831 => std_logic_vector(to_unsigned(21042, 16)), -- 21042 / 0x5232
     832 => std_logic_vector(to_unsigned(37024, 16)), -- 37024 / 0x90a0
     833 => std_logic_vector(to_unsigned(20692, 16)), -- 20692 / 0x50d4 -- last item of row
     834 => std_logic_vector(to_unsigned( 1874, 16)), --  1874 / 0x0752
     835 => std_logic_vector(to_unsigned(40094, 16)), -- 40094 / 0x9c9e
     836 => std_logic_vector(to_unsigned(18704, 16)), -- 18704 / 0x4910
     837 => std_logic_vector(to_unsigned(14474, 16)), -- 14474 / 0x388a
     838 => std_logic_vector(to_unsigned(14004, 16)), -- 14004 / 0x36b4
     839 => std_logic_vector(to_unsigned(11519, 16)), -- 11519 / 0x2cff
     840 => std_logic_vector(to_unsigned(13106, 16)), -- 13106 / 0x3332
     841 => std_logic_vector(to_unsigned(28826, 16)), -- 28826 / 0x709a
     842 => std_logic_vector(to_unsigned(38669, 16)), -- 38669 / 0x970d
     843 => std_logic_vector(to_unsigned(22363, 16)), -- 22363 / 0x575b
     844 => std_logic_vector(to_unsigned(30255, 16)), -- 30255 / 0x762f
     845 => std_logic_vector(to_unsigned(31105, 16)), -- 31105 / 0x7981 -- last item of row
     846 => std_logic_vector(to_unsigned(22254, 16)), -- 22254 / 0x56ee
     847 => std_logic_vector(to_unsigned(40564, 16)), -- 40564 / 0x9e74
     848 => std_logic_vector(to_unsigned(22645, 16)), -- 22645 / 0x5875
     849 => std_logic_vector(to_unsigned(22532, 16)), -- 22532 / 0x5804
     850 => std_logic_vector(to_unsigned( 6134, 16)), --  6134 / 0x17f6
     851 => std_logic_vector(to_unsigned( 9176, 16)), --  9176 / 0x23d8
     852 => std_logic_vector(to_unsigned(39998, 16)), -- 39998 / 0x9c3e
     853 => std_logic_vector(to_unsigned(23892, 16)), -- 23892 / 0x5d54
     854 => std_logic_vector(to_unsigned( 8937, 16)), --  8937 / 0x22e9
     855 => std_logic_vector(to_unsigned(15608, 16)), -- 15608 / 0x3cf8
     856 => std_logic_vector(to_unsigned(16854, 16)), -- 16854 / 0x41d6
     857 => std_logic_vector(to_unsigned(31009, 16)), -- 31009 / 0x7921 -- last item of row
     858 => std_logic_vector(to_unsigned( 8037, 16)), --  8037 / 0x1f65
     859 => std_logic_vector(to_unsigned(40401, 16)), -- 40401 / 0x9dd1
     860 => std_logic_vector(to_unsigned(13550, 16)), -- 13550 / 0x34ee
     861 => std_logic_vector(to_unsigned(19526, 16)), -- 19526 / 0x4c46
     862 => std_logic_vector(to_unsigned(41902, 16)), -- 41902 / 0xa3ae
     863 => std_logic_vector(to_unsigned(28782, 16)), -- 28782 / 0x706e
     864 => std_logic_vector(to_unsigned(13304, 16)), -- 13304 / 0x33f8
     865 => std_logic_vector(to_unsigned(32796, 16)), -- 32796 / 0x801c
     866 => std_logic_vector(to_unsigned(24679, 16)), -- 24679 / 0x6067
     867 => std_logic_vector(to_unsigned(27140, 16)), -- 27140 / 0x6a04
     868 => std_logic_vector(to_unsigned(45980, 16)), -- 45980 / 0xb39c
     869 => std_logic_vector(to_unsigned(10021, 16)), -- 10021 / 0x2725 -- last item of row
     870 => std_logic_vector(to_unsigned(40540, 16)), -- 40540 / 0x9e5c
     871 => std_logic_vector(to_unsigned(44498, 16)), -- 44498 / 0xadd2
     872 => std_logic_vector(to_unsigned(13911, 16)), -- 13911 / 0x3657
     873 => std_logic_vector(to_unsigned(22435, 16)), -- 22435 / 0x57a3
     874 => std_logic_vector(to_unsigned(32701, 16)), -- 32701 / 0x7fbd
     875 => std_logic_vector(to_unsigned(18405, 16)), -- 18405 / 0x47e5
     876 => std_logic_vector(to_unsigned(39929, 16)), -- 39929 / 0x9bf9
     877 => std_logic_vector(to_unsigned(25521, 16)), -- 25521 / 0x63b1
     878 => std_logic_vector(to_unsigned(12497, 16)), -- 12497 / 0x30d1
     879 => std_logic_vector(to_unsigned( 9851, 16)), --  9851 / 0x267b
     880 => std_logic_vector(to_unsigned(39223, 16)), -- 39223 / 0x9937
     881 => std_logic_vector(to_unsigned(34823, 16)), -- 34823 / 0x8807 -- last item of row
     882 => std_logic_vector(to_unsigned(15233, 16)), -- 15233 / 0x3b81
     883 => std_logic_vector(to_unsigned(45333, 16)), -- 45333 / 0xb115
     884 => std_logic_vector(to_unsigned( 5041, 16)), --  5041 / 0x13b1
     885 => std_logic_vector(to_unsigned(44979, 16)), -- 44979 / 0xafb3
     886 => std_logic_vector(to_unsigned(45710, 16)), -- 45710 / 0xb28e
     887 => std_logic_vector(to_unsigned(42150, 16)), -- 42150 / 0xa4a6
     888 => std_logic_vector(to_unsigned(19416, 16)), -- 19416 / 0x4bd8
     889 => std_logic_vector(to_unsigned( 1892, 16)), --  1892 / 0x0764
     890 => std_logic_vector(to_unsigned(23121, 16)), -- 23121 / 0x5a51
     891 => std_logic_vector(to_unsigned(15860, 16)), -- 15860 / 0x3df4
     892 => std_logic_vector(to_unsigned( 8832, 16)), --  8832 / 0x2280
     893 => std_logic_vector(to_unsigned(10308, 16)), -- 10308 / 0x2844 -- last item of row
     894 => std_logic_vector(to_unsigned(10468, 16)), -- 10468 / 0x28e4
     895 => std_logic_vector(to_unsigned(44296, 16)), -- 44296 / 0xad08
     896 => std_logic_vector(to_unsigned( 3611, 16)), --  3611 / 0x0e1b
     897 => std_logic_vector(to_unsigned( 1480, 16)), --  1480 / 0x05c8
     898 => std_logic_vector(to_unsigned(37581, 16)), -- 37581 / 0x92cd
     899 => std_logic_vector(to_unsigned(32254, 16)), -- 32254 / 0x7dfe
     900 => std_logic_vector(to_unsigned(13817, 16)), -- 13817 / 0x35f9
     901 => std_logic_vector(to_unsigned( 6883, 16)), --  6883 / 0x1ae3
     902 => std_logic_vector(to_unsigned(32892, 16)), -- 32892 / 0x807c
     903 => std_logic_vector(to_unsigned(40258, 16)), -- 40258 / 0x9d42
     904 => std_logic_vector(to_unsigned(46538, 16)), -- 46538 / 0xb5ca
     905 => std_logic_vector(to_unsigned(11940, 16)), -- 11940 / 0x2ea4 -- last item of row
     906 => std_logic_vector(to_unsigned( 6705, 16)), --  6705 / 0x1a31
     907 => std_logic_vector(to_unsigned(21634, 16)), -- 21634 / 0x5482
     908 => std_logic_vector(to_unsigned(28150, 16)), -- 28150 / 0x6df6
     909 => std_logic_vector(to_unsigned(43757, 16)), -- 43757 / 0xaaed
     910 => std_logic_vector(to_unsigned(  895, 16)), --   895 / 0x037f
     911 => std_logic_vector(to_unsigned( 6547, 16)), --  6547 / 0x1993
     912 => std_logic_vector(to_unsigned(20970, 16)), -- 20970 / 0x51ea
     913 => std_logic_vector(to_unsigned(28914, 16)), -- 28914 / 0x70f2
     914 => std_logic_vector(to_unsigned(30117, 16)), -- 30117 / 0x75a5
     915 => std_logic_vector(to_unsigned(25736, 16)), -- 25736 / 0x6488
     916 => std_logic_vector(to_unsigned(41734, 16)), -- 41734 / 0xa306
     917 => std_logic_vector(to_unsigned(11392, 16)), -- 11392 / 0x2c80 -- last item of row
     918 => std_logic_vector(to_unsigned(22002, 16)), -- 22002 / 0x55f2
     919 => std_logic_vector(to_unsigned( 5739, 16)), --  5739 / 0x166b
     920 => std_logic_vector(to_unsigned(27210, 16)), -- 27210 / 0x6a4a
     921 => std_logic_vector(to_unsigned(27828, 16)), -- 27828 / 0x6cb4
     922 => std_logic_vector(to_unsigned(34192, 16)), -- 34192 / 0x8590
     923 => std_logic_vector(to_unsigned(37992, 16)), -- 37992 / 0x9468
     924 => std_logic_vector(to_unsigned(10915, 16)), -- 10915 / 0x2aa3
     925 => std_logic_vector(to_unsigned( 6998, 16)), --  6998 / 0x1b56
     926 => std_logic_vector(to_unsigned( 3824, 16)), --  3824 / 0x0ef0
     927 => std_logic_vector(to_unsigned(42130, 16)), -- 42130 / 0xa492
     928 => std_logic_vector(to_unsigned( 4494, 16)), --  4494 / 0x118e
     929 => std_logic_vector(to_unsigned(35739, 16)), -- 35739 / 0x8b9b -- last item of row
     930 => std_logic_vector(to_unsigned( 8515, 16)), --  8515 / 0x2143
     931 => std_logic_vector(to_unsigned( 1191, 16)), --  1191 / 0x04a7
     932 => std_logic_vector(to_unsigned(13642, 16)), -- 13642 / 0x354a
     933 => std_logic_vector(to_unsigned(30950, 16)), -- 30950 / 0x78e6
     934 => std_logic_vector(to_unsigned(25943, 16)), -- 25943 / 0x6557
     935 => std_logic_vector(to_unsigned(12673, 16)), -- 12673 / 0x3181
     936 => std_logic_vector(to_unsigned(16726, 16)), -- 16726 / 0x4156
     937 => std_logic_vector(to_unsigned(34261, 16)), -- 34261 / 0x85d5
     938 => std_logic_vector(to_unsigned(31828, 16)), -- 31828 / 0x7c54
     939 => std_logic_vector(to_unsigned( 3340, 16)), --  3340 / 0x0d0c
     940 => std_logic_vector(to_unsigned( 8747, 16)), --  8747 / 0x222b
     941 => std_logic_vector(to_unsigned(39225, 16)), -- 39225 / 0x9939 -- last item of row
     942 => std_logic_vector(to_unsigned(18979, 16)), -- 18979 / 0x4a23
     943 => std_logic_vector(to_unsigned(17058, 16)), -- 17058 / 0x42a2
     944 => std_logic_vector(to_unsigned(43130, 16)), -- 43130 / 0xa87a
     945 => std_logic_vector(to_unsigned( 4246, 16)), --  4246 / 0x1096
     946 => std_logic_vector(to_unsigned( 4793, 16)), --  4793 / 0x12b9
     947 => std_logic_vector(to_unsigned(44030, 16)), -- 44030 / 0xabfe
     948 => std_logic_vector(to_unsigned(19454, 16)), -- 19454 / 0x4bfe
     949 => std_logic_vector(to_unsigned(29511, 16)), -- 29511 / 0x7347
     950 => std_logic_vector(to_unsigned(47929, 16)), -- 47929 / 0xbb39
     951 => std_logic_vector(to_unsigned(15174, 16)), -- 15174 / 0x3b46
     952 => std_logic_vector(to_unsigned(24333, 16)), -- 24333 / 0x5f0d
     953 => std_logic_vector(to_unsigned(19354, 16)), -- 19354 / 0x4b9a -- last item of row
     954 => std_logic_vector(to_unsigned(16694, 16)), -- 16694 / 0x4136
     955 => std_logic_vector(to_unsigned( 8381, 16)), --  8381 / 0x20bd
     956 => std_logic_vector(to_unsigned(29642, 16)), -- 29642 / 0x73ca
     957 => std_logic_vector(to_unsigned(46516, 16)), -- 46516 / 0xb5b4
     958 => std_logic_vector(to_unsigned(32224, 16)), -- 32224 / 0x7de0
     959 => std_logic_vector(to_unsigned(26344, 16)), -- 26344 / 0x66e8
     960 => std_logic_vector(to_unsigned( 9405, 16)), --  9405 / 0x24bd
     961 => std_logic_vector(to_unsigned(18292, 16)), -- 18292 / 0x4774
     962 => std_logic_vector(to_unsigned(12437, 16)), -- 12437 / 0x3095
     963 => std_logic_vector(to_unsigned(27316, 16)), -- 27316 / 0x6ab4
     964 => std_logic_vector(to_unsigned(35466, 16)), -- 35466 / 0x8a8a
     965 => std_logic_vector(to_unsigned(41992, 16)), -- 41992 / 0xa408 -- last item of row
     966 => std_logic_vector(to_unsigned(15642, 16)), -- 15642 / 0x3d1a
     967 => std_logic_vector(to_unsigned( 5871, 16)), --  5871 / 0x16ef
     968 => std_logic_vector(to_unsigned(46489, 16)), -- 46489 / 0xb599
     969 => std_logic_vector(to_unsigned(26723, 16)), -- 26723 / 0x6863
     970 => std_logic_vector(to_unsigned(23396, 16)), -- 23396 / 0x5b64
     971 => std_logic_vector(to_unsigned( 7257, 16)), --  7257 / 0x1c59
     972 => std_logic_vector(to_unsigned( 8974, 16)), --  8974 / 0x230e
     973 => std_logic_vector(to_unsigned( 3156, 16)), --  3156 / 0x0c54
     974 => std_logic_vector(to_unsigned(37420, 16)), -- 37420 / 0x922c
     975 => std_logic_vector(to_unsigned(44823, 16)), -- 44823 / 0xaf17
     976 => std_logic_vector(to_unsigned(35423, 16)), -- 35423 / 0x8a5f
     977 => std_logic_vector(to_unsigned(13541, 16)), -- 13541 / 0x34e5 -- last item of row
     978 => std_logic_vector(to_unsigned(42858, 16)), -- 42858 / 0xa76a
     979 => std_logic_vector(to_unsigned(32008, 16)), -- 32008 / 0x7d08
     980 => std_logic_vector(to_unsigned(41282, 16)), -- 41282 / 0xa142
     981 => std_logic_vector(to_unsigned(38773, 16)), -- 38773 / 0x9775
     982 => std_logic_vector(to_unsigned(26570, 16)), -- 26570 / 0x67ca
     983 => std_logic_vector(to_unsigned( 2702, 16)), --  2702 / 0x0a8e
     984 => std_logic_vector(to_unsigned(27260, 16)), -- 27260 / 0x6a7c
     985 => std_logic_vector(to_unsigned(46974, 16)), -- 46974 / 0xb77e
     986 => std_logic_vector(to_unsigned( 1469, 16)), --  1469 / 0x05bd
     987 => std_logic_vector(to_unsigned(20887, 16)), -- 20887 / 0x5197
     988 => std_logic_vector(to_unsigned(27426, 16)), -- 27426 / 0x6b22
     989 => std_logic_vector(to_unsigned(38553, 16)), -- 38553 / 0x9699 -- last item of row
     990 => std_logic_vector(to_unsigned(22152, 16)), -- 22152 / 0x5688
     991 => std_logic_vector(to_unsigned(24261, 16)), -- 24261 / 0x5ec5
     992 => std_logic_vector(to_unsigned( 8297, 16)), --  8297 / 0x2069 -- last item of row
     993 => std_logic_vector(to_unsigned(19347, 16)), -- 19347 / 0x4b93
     994 => std_logic_vector(to_unsigned( 9978, 16)), --  9978 / 0x26fa
     995 => std_logic_vector(to_unsigned(27802, 16)), -- 27802 / 0x6c9a -- last item of row
     996 => std_logic_vector(to_unsigned(34991, 16)), -- 34991 / 0x88af
     997 => std_logic_vector(to_unsigned( 6354, 16)), --  6354 / 0x18d2
     998 => std_logic_vector(to_unsigned(33561, 16)), -- 33561 / 0x8319 -- last item of row
     999 => std_logic_vector(to_unsigned(29782, 16)), -- 29782 / 0x7456
    1000 => std_logic_vector(to_unsigned(30875, 16)), -- 30875 / 0x789b
    1001 => std_logic_vector(to_unsigned(29523, 16)), -- 29523 / 0x7353 -- last item of row
    1002 => std_logic_vector(to_unsigned( 9278, 16)), --  9278 / 0x243e
    1003 => std_logic_vector(to_unsigned(48512, 16)), -- 48512 / 0xbd80
    1004 => std_logic_vector(to_unsigned(14349, 16)), -- 14349 / 0x380d -- last item of row
    1005 => std_logic_vector(to_unsigned(38061, 16)), -- 38061 / 0x94ad
    1006 => std_logic_vector(to_unsigned( 4165, 16)), --  4165 / 0x1045
    1007 => std_logic_vector(to_unsigned(43878, 16)), -- 43878 / 0xab66 -- last item of row
    1008 => std_logic_vector(to_unsigned( 8548, 16)), --  8548 / 0x2164
    1009 => std_logic_vector(to_unsigned(33172, 16)), -- 33172 / 0x8194
    1010 => std_logic_vector(to_unsigned(34410, 16)), -- 34410 / 0x866a -- last item of row
    1011 => std_logic_vector(to_unsigned(22535, 16)), -- 22535 / 0x5807
    1012 => std_logic_vector(to_unsigned(28811, 16)), -- 28811 / 0x708b
    1013 => std_logic_vector(to_unsigned(23950, 16)), -- 23950 / 0x5d8e -- last item of row
    1014 => std_logic_vector(to_unsigned(20439, 16)), -- 20439 / 0x4fd7
    1015 => std_logic_vector(to_unsigned( 4027, 16)), --  4027 / 0x0fbb
    1016 => std_logic_vector(to_unsigned(24186, 16)), -- 24186 / 0x5e7a -- last item of row
    1017 => std_logic_vector(to_unsigned(38618, 16)), -- 38618 / 0x96da
    1018 => std_logic_vector(to_unsigned( 8187, 16)), --  8187 / 0x1ffb
    1019 => std_logic_vector(to_unsigned(30947, 16)), -- 30947 / 0x78e3 -- last item of row
    1020 => std_logic_vector(to_unsigned(35538, 16)), -- 35538 / 0x8ad2
    1021 => std_logic_vector(to_unsigned(43880, 16)), -- 43880 / 0xab68
    1022 => std_logic_vector(to_unsigned(21459, 16)), -- 21459 / 0x53d3 -- last item of row
    1023 => std_logic_vector(to_unsigned( 7091, 16)), --  7091 / 0x1bb3
    1024 => std_logic_vector(to_unsigned(45616, 16)), -- 45616 / 0xb230
    1025 => std_logic_vector(to_unsigned(15063, 16)), -- 15063 / 0x3ad7 -- last item of row
    1026 => std_logic_vector(to_unsigned( 5505, 16)), --  5505 / 0x1581
    1027 => std_logic_vector(to_unsigned( 9315, 16)), --  9315 / 0x2463
    1028 => std_logic_vector(to_unsigned(21908, 16)), -- 21908 / 0x5594 -- last item of row
    1029 => std_logic_vector(to_unsigned(36046, 16)), -- 36046 / 0x8cce
    1030 => std_logic_vector(to_unsigned(32914, 16)), -- 32914 / 0x8092
    1031 => std_logic_vector(to_unsigned(11836, 16)), -- 11836 / 0x2e3c -- last item of row
    1032 => std_logic_vector(to_unsigned( 7304, 16)), --  7304 / 0x1c88
    1033 => std_logic_vector(to_unsigned(39782, 16)), -- 39782 / 0x9b66
    1034 => std_logic_vector(to_unsigned(33721, 16)), -- 33721 / 0x83b9 -- last item of row
    1035 => std_logic_vector(to_unsigned(16905, 16)), -- 16905 / 0x4209
    1036 => std_logic_vector(to_unsigned(29962, 16)), -- 29962 / 0x750a
    1037 => std_logic_vector(to_unsigned(12980, 16)), -- 12980 / 0x32b4 -- last item of row
    1038 => std_logic_vector(to_unsigned(11171, 16)), -- 11171 / 0x2ba3
    1039 => std_logic_vector(to_unsigned(23709, 16)), -- 23709 / 0x5c9d
    1040 => std_logic_vector(to_unsigned(22460, 16)), -- 22460 / 0x57bc -- last item of row
    1041 => std_logic_vector(to_unsigned(34541, 16)), -- 34541 / 0x86ed
    1042 => std_logic_vector(to_unsigned( 9937, 16)), --  9937 / 0x26d1
    1043 => std_logic_vector(to_unsigned(44500, 16)), -- 44500 / 0xadd4 -- last item of row
    1044 => std_logic_vector(to_unsigned(14035, 16)), -- 14035 / 0x36d3
    1045 => std_logic_vector(to_unsigned(47316, 16)), -- 47316 / 0xb8d4
    1046 => std_logic_vector(to_unsigned( 8815, 16)), --  8815 / 0x226f -- last item of row
    1047 => std_logic_vector(to_unsigned(15057, 16)), -- 15057 / 0x3ad1
    1048 => std_logic_vector(to_unsigned(45482, 16)), -- 45482 / 0xb1aa
    1049 => std_logic_vector(to_unsigned(24461, 16)), -- 24461 / 0x5f8d -- last item of row
    1050 => std_logic_vector(to_unsigned(30518, 16)), -- 30518 / 0x7736
    1051 => std_logic_vector(to_unsigned(36877, 16)), -- 36877 / 0x900d
    1052 => std_logic_vector(to_unsigned(  879, 16)), --   879 / 0x036f -- last item of row
    1053 => std_logic_vector(to_unsigned( 7583, 16)), --  7583 / 0x1d9f
    1054 => std_logic_vector(to_unsigned(13364, 16)), -- 13364 / 0x3434
    1055 => std_logic_vector(to_unsigned(24332, 16)), -- 24332 / 0x5f0c -- last item of row
    1056 => std_logic_vector(to_unsigned(  448, 16)), --   448 / 0x01c0
    1057 => std_logic_vector(to_unsigned(27056, 16)), -- 27056 / 0x69b0
    1058 => std_logic_vector(to_unsigned( 4682, 16)), --  4682 / 0x124a -- last item of row
    1059 => std_logic_vector(to_unsigned(12083, 16)), -- 12083 / 0x2f33
    1060 => std_logic_vector(to_unsigned(31378, 16)), -- 31378 / 0x7a92
    1061 => std_logic_vector(to_unsigned(21670, 16)), -- 21670 / 0x54a6 -- last item of row
    1062 => std_logic_vector(to_unsigned( 1159, 16)), --  1159 / 0x0487
    1063 => std_logic_vector(to_unsigned(18031, 16)), -- 18031 / 0x466f
    1064 => std_logic_vector(to_unsigned( 2221, 16)), --  2221 / 0x08ad -- last item of row
    1065 => std_logic_vector(to_unsigned(17028, 16)), -- 17028 / 0x4284
    1066 => std_logic_vector(to_unsigned(38715, 16)), -- 38715 / 0x973b
    1067 => std_logic_vector(to_unsigned( 9350, 16)), --  9350 / 0x2486 -- last item of row
    1068 => std_logic_vector(to_unsigned(17343, 16)), -- 17343 / 0x43bf
    1069 => std_logic_vector(to_unsigned(24530, 16)), -- 24530 / 0x5fd2
    1070 => std_logic_vector(to_unsigned(29574, 16)), -- 29574 / 0x7386 -- last item of row
    1071 => std_logic_vector(to_unsigned(46128, 16)), -- 46128 / 0xb430
    1072 => std_logic_vector(to_unsigned(31039, 16)), -- 31039 / 0x793f
    1073 => std_logic_vector(to_unsigned(32818, 16)), -- 32818 / 0x8032 -- last item of row
    1074 => std_logic_vector(to_unsigned(20373, 16)), -- 20373 / 0x4f95
    1075 => std_logic_vector(to_unsigned(36967, 16)), -- 36967 / 0x9067
    1076 => std_logic_vector(to_unsigned(18345, 16)), -- 18345 / 0x47a9 -- last item of row
    1077 => std_logic_vector(to_unsigned(46685, 16)), -- 46685 / 0xb65d
    1078 => std_logic_vector(to_unsigned(20622, 16)), -- 20622 / 0x508e
    1079 => std_logic_vector(to_unsigned(32806, 16)), -- 32806 / 0x8026 -- last item of row
    -- Table for fecframe_normal, C2_3
    1080 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    1081 => std_logic_vector(to_unsigned(10491, 16)), -- 10491 / 0x28fb
    1082 => std_logic_vector(to_unsigned(16043, 16)), -- 16043 / 0x3eab
    1083 => std_logic_vector(to_unsigned(  506, 16)), --   506 / 0x01fa
    1084 => std_logic_vector(to_unsigned(12826, 16)), -- 12826 / 0x321a
    1085 => std_logic_vector(to_unsigned( 8065, 16)), --  8065 / 0x1f81
    1086 => std_logic_vector(to_unsigned( 8226, 16)), --  8226 / 0x2022
    1087 => std_logic_vector(to_unsigned( 2767, 16)), --  2767 / 0x0acf
    1088 => std_logic_vector(to_unsigned(  240, 16)), --   240 / 0x00f0
    1089 => std_logic_vector(to_unsigned(18673, 16)), -- 18673 / 0x48f1
    1090 => std_logic_vector(to_unsigned( 9279, 16)), --  9279 / 0x243f
    1091 => std_logic_vector(to_unsigned(10579, 16)), -- 10579 / 0x2953
    1092 => std_logic_vector(to_unsigned(20928, 16)), -- 20928 / 0x51c0 -- last item of row
    1093 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    1094 => std_logic_vector(to_unsigned(17819, 16)), -- 17819 / 0x459b
    1095 => std_logic_vector(to_unsigned( 8313, 16)), --  8313 / 0x2079
    1096 => std_logic_vector(to_unsigned( 6433, 16)), --  6433 / 0x1921
    1097 => std_logic_vector(to_unsigned( 6224, 16)), --  6224 / 0x1850
    1098 => std_logic_vector(to_unsigned( 5120, 16)), --  5120 / 0x1400
    1099 => std_logic_vector(to_unsigned( 5824, 16)), --  5824 / 0x16c0
    1100 => std_logic_vector(to_unsigned(12812, 16)), -- 12812 / 0x320c
    1101 => std_logic_vector(to_unsigned(17187, 16)), -- 17187 / 0x4323
    1102 => std_logic_vector(to_unsigned( 9940, 16)), --  9940 / 0x26d4
    1103 => std_logic_vector(to_unsigned(13447, 16)), -- 13447 / 0x3487
    1104 => std_logic_vector(to_unsigned(13825, 16)), -- 13825 / 0x3601
    1105 => std_logic_vector(to_unsigned(18483, 16)), -- 18483 / 0x4833 -- last item of row
    1106 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    1107 => std_logic_vector(to_unsigned(17957, 16)), -- 17957 / 0x4625
    1108 => std_logic_vector(to_unsigned( 6024, 16)), --  6024 / 0x1788
    1109 => std_logic_vector(to_unsigned( 8681, 16)), --  8681 / 0x21e9
    1110 => std_logic_vector(to_unsigned(18628, 16)), -- 18628 / 0x48c4
    1111 => std_logic_vector(to_unsigned(12794, 16)), -- 12794 / 0x31fa
    1112 => std_logic_vector(to_unsigned( 5915, 16)), --  5915 / 0x171b
    1113 => std_logic_vector(to_unsigned(14576, 16)), -- 14576 / 0x38f0
    1114 => std_logic_vector(to_unsigned(10970, 16)), -- 10970 / 0x2ada
    1115 => std_logic_vector(to_unsigned(12064, 16)), -- 12064 / 0x2f20
    1116 => std_logic_vector(to_unsigned(20437, 16)), -- 20437 / 0x4fd5
    1117 => std_logic_vector(to_unsigned( 4455, 16)), --  4455 / 0x1167
    1118 => std_logic_vector(to_unsigned( 7151, 16)), --  7151 / 0x1bef -- last item of row
    1119 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    1120 => std_logic_vector(to_unsigned(19777, 16)), -- 19777 / 0x4d41
    1121 => std_logic_vector(to_unsigned( 6183, 16)), --  6183 / 0x1827
    1122 => std_logic_vector(to_unsigned( 9972, 16)), --  9972 / 0x26f4
    1123 => std_logic_vector(to_unsigned(14536, 16)), -- 14536 / 0x38c8
    1124 => std_logic_vector(to_unsigned( 8182, 16)), --  8182 / 0x1ff6
    1125 => std_logic_vector(to_unsigned(17749, 16)), -- 17749 / 0x4555
    1126 => std_logic_vector(to_unsigned(11341, 16)), -- 11341 / 0x2c4d
    1127 => std_logic_vector(to_unsigned( 5556, 16)), --  5556 / 0x15b4
    1128 => std_logic_vector(to_unsigned( 4379, 16)), --  4379 / 0x111b
    1129 => std_logic_vector(to_unsigned(17434, 16)), -- 17434 / 0x441a
    1130 => std_logic_vector(to_unsigned(15477, 16)), -- 15477 / 0x3c75
    1131 => std_logic_vector(to_unsigned(18532, 16)), -- 18532 / 0x4864 -- last item of row
    1132 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    1133 => std_logic_vector(to_unsigned( 4651, 16)), --  4651 / 0x122b
    1134 => std_logic_vector(to_unsigned(19689, 16)), -- 19689 / 0x4ce9
    1135 => std_logic_vector(to_unsigned( 1608, 16)), --  1608 / 0x0648
    1136 => std_logic_vector(to_unsigned(  659, 16)), --   659 / 0x0293
    1137 => std_logic_vector(to_unsigned(16707, 16)), -- 16707 / 0x4143
    1138 => std_logic_vector(to_unsigned(14335, 16)), -- 14335 / 0x37ff
    1139 => std_logic_vector(to_unsigned( 6143, 16)), --  6143 / 0x17ff
    1140 => std_logic_vector(to_unsigned( 3058, 16)), --  3058 / 0x0bf2
    1141 => std_logic_vector(to_unsigned(14618, 16)), -- 14618 / 0x391a
    1142 => std_logic_vector(to_unsigned(17894, 16)), -- 17894 / 0x45e6
    1143 => std_logic_vector(to_unsigned(20684, 16)), -- 20684 / 0x50cc
    1144 => std_logic_vector(to_unsigned( 5306, 16)), --  5306 / 0x14ba -- last item of row
    1145 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    1146 => std_logic_vector(to_unsigned( 9778, 16)), --  9778 / 0x2632
    1147 => std_logic_vector(to_unsigned( 2552, 16)), --  2552 / 0x09f8
    1148 => std_logic_vector(to_unsigned(12096, 16)), -- 12096 / 0x2f40
    1149 => std_logic_vector(to_unsigned(12369, 16)), -- 12369 / 0x3051
    1150 => std_logic_vector(to_unsigned(15198, 16)), -- 15198 / 0x3b5e
    1151 => std_logic_vector(to_unsigned(16890, 16)), -- 16890 / 0x41fa
    1152 => std_logic_vector(to_unsigned( 4851, 16)), --  4851 / 0x12f3
    1153 => std_logic_vector(to_unsigned( 3109, 16)), --  3109 / 0x0c25
    1154 => std_logic_vector(to_unsigned( 1700, 16)), --  1700 / 0x06a4
    1155 => std_logic_vector(to_unsigned(18725, 16)), -- 18725 / 0x4925
    1156 => std_logic_vector(to_unsigned( 1997, 16)), --  1997 / 0x07cd
    1157 => std_logic_vector(to_unsigned(15882, 16)), -- 15882 / 0x3e0a -- last item of row
    1158 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    1159 => std_logic_vector(to_unsigned(  486, 16)), --   486 / 0x01e6
    1160 => std_logic_vector(to_unsigned( 6111, 16)), --  6111 / 0x17df
    1161 => std_logic_vector(to_unsigned(13743, 16)), -- 13743 / 0x35af
    1162 => std_logic_vector(to_unsigned(11537, 16)), -- 11537 / 0x2d11
    1163 => std_logic_vector(to_unsigned( 5591, 16)), --  5591 / 0x15d7
    1164 => std_logic_vector(to_unsigned( 7433, 16)), --  7433 / 0x1d09
    1165 => std_logic_vector(to_unsigned(15227, 16)), -- 15227 / 0x3b7b
    1166 => std_logic_vector(to_unsigned(14145, 16)), -- 14145 / 0x3741
    1167 => std_logic_vector(to_unsigned( 1483, 16)), --  1483 / 0x05cb
    1168 => std_logic_vector(to_unsigned( 3887, 16)), --  3887 / 0x0f2f
    1169 => std_logic_vector(to_unsigned(17431, 16)), -- 17431 / 0x4417
    1170 => std_logic_vector(to_unsigned(12430, 16)), -- 12430 / 0x308e -- last item of row
    1171 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    1172 => std_logic_vector(to_unsigned(20647, 16)), -- 20647 / 0x50a7
    1173 => std_logic_vector(to_unsigned(14311, 16)), -- 14311 / 0x37e7
    1174 => std_logic_vector(to_unsigned(11734, 16)), -- 11734 / 0x2dd6
    1175 => std_logic_vector(to_unsigned( 4180, 16)), --  4180 / 0x1054
    1176 => std_logic_vector(to_unsigned( 8110, 16)), --  8110 / 0x1fae
    1177 => std_logic_vector(to_unsigned( 5525, 16)), --  5525 / 0x1595
    1178 => std_logic_vector(to_unsigned(12141, 16)), -- 12141 / 0x2f6d
    1179 => std_logic_vector(to_unsigned(15761, 16)), -- 15761 / 0x3d91
    1180 => std_logic_vector(to_unsigned(18661, 16)), -- 18661 / 0x48e5
    1181 => std_logic_vector(to_unsigned(18441, 16)), -- 18441 / 0x4809
    1182 => std_logic_vector(to_unsigned(10569, 16)), -- 10569 / 0x2949
    1183 => std_logic_vector(to_unsigned( 8192, 16)), --  8192 / 0x2000 -- last item of row
    1184 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    1185 => std_logic_vector(to_unsigned( 3791, 16)), --  3791 / 0x0ecf
    1186 => std_logic_vector(to_unsigned(14759, 16)), -- 14759 / 0x39a7
    1187 => std_logic_vector(to_unsigned(15264, 16)), -- 15264 / 0x3ba0
    1188 => std_logic_vector(to_unsigned(19918, 16)), -- 19918 / 0x4dce
    1189 => std_logic_vector(to_unsigned(10132, 16)), -- 10132 / 0x2794
    1190 => std_logic_vector(to_unsigned( 9062, 16)), --  9062 / 0x2366
    1191 => std_logic_vector(to_unsigned(10010, 16)), -- 10010 / 0x271a
    1192 => std_logic_vector(to_unsigned(12786, 16)), -- 12786 / 0x31f2
    1193 => std_logic_vector(to_unsigned(10675, 16)), -- 10675 / 0x29b3
    1194 => std_logic_vector(to_unsigned( 9682, 16)), --  9682 / 0x25d2
    1195 => std_logic_vector(to_unsigned(19246, 16)), -- 19246 / 0x4b2e
    1196 => std_logic_vector(to_unsigned( 5454, 16)), --  5454 / 0x154e -- last item of row
    1197 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    1198 => std_logic_vector(to_unsigned(19525, 16)), -- 19525 / 0x4c45
    1199 => std_logic_vector(to_unsigned( 9485, 16)), --  9485 / 0x250d
    1200 => std_logic_vector(to_unsigned( 7777, 16)), --  7777 / 0x1e61
    1201 => std_logic_vector(to_unsigned(19999, 16)), -- 19999 / 0x4e1f
    1202 => std_logic_vector(to_unsigned( 8378, 16)), --  8378 / 0x20ba
    1203 => std_logic_vector(to_unsigned( 9209, 16)), --  9209 / 0x23f9
    1204 => std_logic_vector(to_unsigned( 3163, 16)), --  3163 / 0x0c5b
    1205 => std_logic_vector(to_unsigned(20232, 16)), -- 20232 / 0x4f08
    1206 => std_logic_vector(to_unsigned( 6690, 16)), --  6690 / 0x1a22
    1207 => std_logic_vector(to_unsigned(16518, 16)), -- 16518 / 0x4086
    1208 => std_logic_vector(to_unsigned(  716, 16)), --   716 / 0x02cc
    1209 => std_logic_vector(to_unsigned( 7353, 16)), --  7353 / 0x1cb9 -- last item of row
    1210 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    1211 => std_logic_vector(to_unsigned( 4588, 16)), --  4588 / 0x11ec
    1212 => std_logic_vector(to_unsigned( 6709, 16)), --  6709 / 0x1a35
    1213 => std_logic_vector(to_unsigned(20202, 16)), -- 20202 / 0x4eea
    1214 => std_logic_vector(to_unsigned(10905, 16)), -- 10905 / 0x2a99
    1215 => std_logic_vector(to_unsigned(  915, 16)), --   915 / 0x0393
    1216 => std_logic_vector(to_unsigned( 4317, 16)), --  4317 / 0x10dd
    1217 => std_logic_vector(to_unsigned(11073, 16)), -- 11073 / 0x2b41
    1218 => std_logic_vector(to_unsigned(13576, 16)), -- 13576 / 0x3508
    1219 => std_logic_vector(to_unsigned(16433, 16)), -- 16433 / 0x4031
    1220 => std_logic_vector(to_unsigned(  368, 16)), --   368 / 0x0170
    1221 => std_logic_vector(to_unsigned( 3508, 16)), --  3508 / 0x0db4
    1222 => std_logic_vector(to_unsigned(21171, 16)), -- 21171 / 0x52b3 -- last item of row
    1223 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    1224 => std_logic_vector(to_unsigned(14072, 16)), -- 14072 / 0x36f8
    1225 => std_logic_vector(to_unsigned( 4033, 16)), --  4033 / 0x0fc1
    1226 => std_logic_vector(to_unsigned(19959, 16)), -- 19959 / 0x4df7
    1227 => std_logic_vector(to_unsigned(12608, 16)), -- 12608 / 0x3140
    1228 => std_logic_vector(to_unsigned(  631, 16)), --   631 / 0x0277
    1229 => std_logic_vector(to_unsigned(19494, 16)), -- 19494 / 0x4c26
    1230 => std_logic_vector(to_unsigned(14160, 16)), -- 14160 / 0x3750
    1231 => std_logic_vector(to_unsigned( 8249, 16)), --  8249 / 0x2039
    1232 => std_logic_vector(to_unsigned(10223, 16)), -- 10223 / 0x27ef
    1233 => std_logic_vector(to_unsigned(21504, 16)), -- 21504 / 0x5400
    1234 => std_logic_vector(to_unsigned(12395, 16)), -- 12395 / 0x306b
    1235 => std_logic_vector(to_unsigned( 4322, 16)), --  4322 / 0x10e2 -- last item of row
    1236 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    1237 => std_logic_vector(to_unsigned(13800, 16)), -- 13800 / 0x35e8
    1238 => std_logic_vector(to_unsigned(14161, 16)), -- 14161 / 0x3751 -- last item of row
    1239 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    1240 => std_logic_vector(to_unsigned( 2948, 16)), --  2948 / 0x0b84
    1241 => std_logic_vector(to_unsigned( 9647, 16)), --  9647 / 0x25af -- last item of row
    1242 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    1243 => std_logic_vector(to_unsigned(14693, 16)), -- 14693 / 0x3965
    1244 => std_logic_vector(to_unsigned(16027, 16)), -- 16027 / 0x3e9b -- last item of row
    1245 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    1246 => std_logic_vector(to_unsigned(20506, 16)), -- 20506 / 0x501a
    1247 => std_logic_vector(to_unsigned(11082, 16)), -- 11082 / 0x2b4a -- last item of row
    1248 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    1249 => std_logic_vector(to_unsigned( 1143, 16)), --  1143 / 0x0477
    1250 => std_logic_vector(to_unsigned( 9020, 16)), --  9020 / 0x233c -- last item of row
    1251 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    1252 => std_logic_vector(to_unsigned(13501, 16)), -- 13501 / 0x34bd
    1253 => std_logic_vector(to_unsigned( 4014, 16)), --  4014 / 0x0fae -- last item of row
    1254 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    1255 => std_logic_vector(to_unsigned( 1548, 16)), --  1548 / 0x060c
    1256 => std_logic_vector(to_unsigned( 2190, 16)), --  2190 / 0x088e -- last item of row
    1257 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    1258 => std_logic_vector(to_unsigned(12216, 16)), -- 12216 / 0x2fb8
    1259 => std_logic_vector(to_unsigned(21556, 16)), -- 21556 / 0x5434 -- last item of row
    1260 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    1261 => std_logic_vector(to_unsigned( 2095, 16)), --  2095 / 0x082f
    1262 => std_logic_vector(to_unsigned(19897, 16)), -- 19897 / 0x4db9 -- last item of row
    1263 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    1264 => std_logic_vector(to_unsigned( 4189, 16)), --  4189 / 0x105d
    1265 => std_logic_vector(to_unsigned( 7958, 16)), --  7958 / 0x1f16 -- last item of row
    1266 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    1267 => std_logic_vector(to_unsigned(15940, 16)), -- 15940 / 0x3e44
    1268 => std_logic_vector(to_unsigned(10048, 16)), -- 10048 / 0x2740 -- last item of row
    1269 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    1270 => std_logic_vector(to_unsigned(  515, 16)), --   515 / 0x0203
    1271 => std_logic_vector(to_unsigned(12614, 16)), -- 12614 / 0x3146 -- last item of row
    1272 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    1273 => std_logic_vector(to_unsigned( 8501, 16)), --  8501 / 0x2135
    1274 => std_logic_vector(to_unsigned( 8450, 16)), --  8450 / 0x2102 -- last item of row
    1275 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    1276 => std_logic_vector(to_unsigned(17595, 16)), -- 17595 / 0x44bb
    1277 => std_logic_vector(to_unsigned(16784, 16)), -- 16784 / 0x4190 -- last item of row
    1278 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    1279 => std_logic_vector(to_unsigned( 5913, 16)), --  5913 / 0x1719
    1280 => std_logic_vector(to_unsigned( 8495, 16)), --  8495 / 0x212f -- last item of row
    1281 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    1282 => std_logic_vector(to_unsigned(16394, 16)), -- 16394 / 0x400a
    1283 => std_logic_vector(to_unsigned(10423, 16)), -- 10423 / 0x28b7 -- last item of row
    1284 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    1285 => std_logic_vector(to_unsigned( 7409, 16)), --  7409 / 0x1cf1
    1286 => std_logic_vector(to_unsigned( 6981, 16)), --  6981 / 0x1b45 -- last item of row
    1287 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    1288 => std_logic_vector(to_unsigned( 6678, 16)), --  6678 / 0x1a16
    1289 => std_logic_vector(to_unsigned(15939, 16)), -- 15939 / 0x3e43 -- last item of row
    1290 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    1291 => std_logic_vector(to_unsigned(20344, 16)), -- 20344 / 0x4f78
    1292 => std_logic_vector(to_unsigned(12987, 16)), -- 12987 / 0x32bb -- last item of row
    1293 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    1294 => std_logic_vector(to_unsigned( 2510, 16)), --  2510 / 0x09ce
    1295 => std_logic_vector(to_unsigned(14588, 16)), -- 14588 / 0x38fc -- last item of row
    1296 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    1297 => std_logic_vector(to_unsigned(17918, 16)), -- 17918 / 0x45fe
    1298 => std_logic_vector(to_unsigned( 6655, 16)), --  6655 / 0x19ff -- last item of row
    1299 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    1300 => std_logic_vector(to_unsigned( 6703, 16)), --  6703 / 0x1a2f
    1301 => std_logic_vector(to_unsigned(19451, 16)), -- 19451 / 0x4bfb -- last item of row
    1302 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    1303 => std_logic_vector(to_unsigned(  496, 16)), --   496 / 0x01f0
    1304 => std_logic_vector(to_unsigned( 4217, 16)), --  4217 / 0x1079 -- last item of row
    1305 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    1306 => std_logic_vector(to_unsigned( 7290, 16)), --  7290 / 0x1c7a
    1307 => std_logic_vector(to_unsigned( 5766, 16)), --  5766 / 0x1686 -- last item of row
    1308 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    1309 => std_logic_vector(to_unsigned(10521, 16)), -- 10521 / 0x2919
    1310 => std_logic_vector(to_unsigned( 8925, 16)), --  8925 / 0x22dd -- last item of row
    1311 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    1312 => std_logic_vector(to_unsigned(20379, 16)), -- 20379 / 0x4f9b
    1313 => std_logic_vector(to_unsigned(11905, 16)), -- 11905 / 0x2e81 -- last item of row
    1314 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    1315 => std_logic_vector(to_unsigned( 4090, 16)), --  4090 / 0x0ffa
    1316 => std_logic_vector(to_unsigned( 5838, 16)), --  5838 / 0x16ce -- last item of row
    1317 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    1318 => std_logic_vector(to_unsigned(19082, 16)), -- 19082 / 0x4a8a
    1319 => std_logic_vector(to_unsigned(17040, 16)), -- 17040 / 0x4290 -- last item of row
    1320 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    1321 => std_logic_vector(to_unsigned(20233, 16)), -- 20233 / 0x4f09
    1322 => std_logic_vector(to_unsigned(12352, 16)), -- 12352 / 0x3040 -- last item of row
    1323 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    1324 => std_logic_vector(to_unsigned(19365, 16)), -- 19365 / 0x4ba5
    1325 => std_logic_vector(to_unsigned(19546, 16)), -- 19546 / 0x4c5a -- last item of row
    1326 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    1327 => std_logic_vector(to_unsigned( 6249, 16)), --  6249 / 0x1869
    1328 => std_logic_vector(to_unsigned(19030, 16)), -- 19030 / 0x4a56 -- last item of row
    1329 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    1330 => std_logic_vector(to_unsigned(11037, 16)), -- 11037 / 0x2b1d
    1331 => std_logic_vector(to_unsigned(19193, 16)), -- 19193 / 0x4af9 -- last item of row
    1332 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    1333 => std_logic_vector(to_unsigned(19760, 16)), -- 19760 / 0x4d30
    1334 => std_logic_vector(to_unsigned(11772, 16)), -- 11772 / 0x2dfc -- last item of row
    1335 => std_logic_vector(to_unsigned(   45, 16)), --    45 / 0x002d
    1336 => std_logic_vector(to_unsigned(19644, 16)), -- 19644 / 0x4cbc
    1337 => std_logic_vector(to_unsigned( 7428, 16)), --  7428 / 0x1d04 -- last item of row
    1338 => std_logic_vector(to_unsigned(   46, 16)), --    46 / 0x002e
    1339 => std_logic_vector(to_unsigned(16076, 16)), -- 16076 / 0x3ecc
    1340 => std_logic_vector(to_unsigned( 3521, 16)), --  3521 / 0x0dc1 -- last item of row
    1341 => std_logic_vector(to_unsigned(   47, 16)), --    47 / 0x002f
    1342 => std_logic_vector(to_unsigned(11779, 16)), -- 11779 / 0x2e03
    1343 => std_logic_vector(to_unsigned(21062, 16)), -- 21062 / 0x5246 -- last item of row
    1344 => std_logic_vector(to_unsigned(   48, 16)), --    48 / 0x0030
    1345 => std_logic_vector(to_unsigned(13062, 16)), -- 13062 / 0x3306
    1346 => std_logic_vector(to_unsigned( 9682, 16)), --  9682 / 0x25d2 -- last item of row
    1347 => std_logic_vector(to_unsigned(   49, 16)), --    49 / 0x0031
    1348 => std_logic_vector(to_unsigned( 8934, 16)), --  8934 / 0x22e6
    1349 => std_logic_vector(to_unsigned( 5217, 16)), --  5217 / 0x1461 -- last item of row
    1350 => std_logic_vector(to_unsigned(   50, 16)), --    50 / 0x0032
    1351 => std_logic_vector(to_unsigned(11087, 16)), -- 11087 / 0x2b4f
    1352 => std_logic_vector(to_unsigned( 3319, 16)), --  3319 / 0x0cf7 -- last item of row
    1353 => std_logic_vector(to_unsigned(   51, 16)), --    51 / 0x0033
    1354 => std_logic_vector(to_unsigned(18892, 16)), -- 18892 / 0x49cc
    1355 => std_logic_vector(to_unsigned( 4356, 16)), --  4356 / 0x1104 -- last item of row
    1356 => std_logic_vector(to_unsigned(   52, 16)), --    52 / 0x0034
    1357 => std_logic_vector(to_unsigned( 7894, 16)), --  7894 / 0x1ed6
    1358 => std_logic_vector(to_unsigned( 3898, 16)), --  3898 / 0x0f3a -- last item of row
    1359 => std_logic_vector(to_unsigned(   53, 16)), --    53 / 0x0035
    1360 => std_logic_vector(to_unsigned( 5963, 16)), --  5963 / 0x174b
    1361 => std_logic_vector(to_unsigned( 4360, 16)), --  4360 / 0x1108 -- last item of row
    1362 => std_logic_vector(to_unsigned(   54, 16)), --    54 / 0x0036
    1363 => std_logic_vector(to_unsigned( 7346, 16)), --  7346 / 0x1cb2
    1364 => std_logic_vector(to_unsigned(11726, 16)), -- 11726 / 0x2dce -- last item of row
    1365 => std_logic_vector(to_unsigned(   55, 16)), --    55 / 0x0037
    1366 => std_logic_vector(to_unsigned( 5182, 16)), --  5182 / 0x143e
    1367 => std_logic_vector(to_unsigned( 5609, 16)), --  5609 / 0x15e9 -- last item of row
    1368 => std_logic_vector(to_unsigned(   56, 16)), --    56 / 0x0038
    1369 => std_logic_vector(to_unsigned( 2412, 16)), --  2412 / 0x096c
    1370 => std_logic_vector(to_unsigned(17295, 16)), -- 17295 / 0x438f -- last item of row
    1371 => std_logic_vector(to_unsigned(   57, 16)), --    57 / 0x0039
    1372 => std_logic_vector(to_unsigned( 9845, 16)), --  9845 / 0x2675
    1373 => std_logic_vector(to_unsigned(20494, 16)), -- 20494 / 0x500e -- last item of row
    1374 => std_logic_vector(to_unsigned(   58, 16)), --    58 / 0x003a
    1375 => std_logic_vector(to_unsigned( 6687, 16)), --  6687 / 0x1a1f
    1376 => std_logic_vector(to_unsigned( 1864, 16)), --  1864 / 0x0748 -- last item of row
    1377 => std_logic_vector(to_unsigned(   59, 16)), --    59 / 0x003b
    1378 => std_logic_vector(to_unsigned(20564, 16)), -- 20564 / 0x5054
    1379 => std_logic_vector(to_unsigned( 5216, 16)), --  5216 / 0x1460 -- last item of row
    1380 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    1381 => std_logic_vector(to_unsigned(18226, 16)), -- 18226 / 0x4732
    1382 => std_logic_vector(to_unsigned(17207, 16)), -- 17207 / 0x4337 -- last item of row
    1383 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    1384 => std_logic_vector(to_unsigned( 9380, 16)), --  9380 / 0x24a4
    1385 => std_logic_vector(to_unsigned( 8266, 16)), --  8266 / 0x204a -- last item of row
    1386 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    1387 => std_logic_vector(to_unsigned( 7073, 16)), --  7073 / 0x1ba1
    1388 => std_logic_vector(to_unsigned( 3065, 16)), --  3065 / 0x0bf9 -- last item of row
    1389 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    1390 => std_logic_vector(to_unsigned(18252, 16)), -- 18252 / 0x474c
    1391 => std_logic_vector(to_unsigned(13437, 16)), -- 13437 / 0x347d -- last item of row
    1392 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    1393 => std_logic_vector(to_unsigned( 9161, 16)), --  9161 / 0x23c9
    1394 => std_logic_vector(to_unsigned(15642, 16)), -- 15642 / 0x3d1a -- last item of row
    1395 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    1396 => std_logic_vector(to_unsigned(10714, 16)), -- 10714 / 0x29da
    1397 => std_logic_vector(to_unsigned(10153, 16)), -- 10153 / 0x27a9 -- last item of row
    1398 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    1399 => std_logic_vector(to_unsigned(11585, 16)), -- 11585 / 0x2d41
    1400 => std_logic_vector(to_unsigned( 9078, 16)), --  9078 / 0x2376 -- last item of row
    1401 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    1402 => std_logic_vector(to_unsigned( 5359, 16)), --  5359 / 0x14ef
    1403 => std_logic_vector(to_unsigned( 9418, 16)), --  9418 / 0x24ca -- last item of row
    1404 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    1405 => std_logic_vector(to_unsigned( 9024, 16)), --  9024 / 0x2340
    1406 => std_logic_vector(to_unsigned( 9515, 16)), --  9515 / 0x252b -- last item of row
    1407 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    1408 => std_logic_vector(to_unsigned( 1206, 16)), --  1206 / 0x04b6
    1409 => std_logic_vector(to_unsigned(16354, 16)), -- 16354 / 0x3fe2 -- last item of row
    1410 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    1411 => std_logic_vector(to_unsigned(14994, 16)), -- 14994 / 0x3a92
    1412 => std_logic_vector(to_unsigned( 1102, 16)), --  1102 / 0x044e -- last item of row
    1413 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    1414 => std_logic_vector(to_unsigned( 9375, 16)), --  9375 / 0x249f
    1415 => std_logic_vector(to_unsigned(20796, 16)), -- 20796 / 0x513c -- last item of row
    1416 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    1417 => std_logic_vector(to_unsigned(15964, 16)), -- 15964 / 0x3e5c
    1418 => std_logic_vector(to_unsigned( 6027, 16)), --  6027 / 0x178b -- last item of row
    1419 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    1420 => std_logic_vector(to_unsigned(14789, 16)), -- 14789 / 0x39c5
    1421 => std_logic_vector(to_unsigned( 6452, 16)), --  6452 / 0x1934 -- last item of row
    1422 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    1423 => std_logic_vector(to_unsigned( 8002, 16)), --  8002 / 0x1f42
    1424 => std_logic_vector(to_unsigned(18591, 16)), -- 18591 / 0x489f -- last item of row
    1425 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    1426 => std_logic_vector(to_unsigned(14742, 16)), -- 14742 / 0x3996
    1427 => std_logic_vector(to_unsigned(14089, 16)), -- 14089 / 0x3709 -- last item of row
    1428 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    1429 => std_logic_vector(to_unsigned(  253, 16)), --   253 / 0x00fd
    1430 => std_logic_vector(to_unsigned( 3045, 16)), --  3045 / 0x0be5 -- last item of row
    1431 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    1432 => std_logic_vector(to_unsigned( 1274, 16)), --  1274 / 0x04fa
    1433 => std_logic_vector(to_unsigned(19286, 16)), -- 19286 / 0x4b56 -- last item of row
    1434 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    1435 => std_logic_vector(to_unsigned(14777, 16)), -- 14777 / 0x39b9
    1436 => std_logic_vector(to_unsigned( 2044, 16)), --  2044 / 0x07fc -- last item of row
    1437 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    1438 => std_logic_vector(to_unsigned(13920, 16)), -- 13920 / 0x3660
    1439 => std_logic_vector(to_unsigned( 9900, 16)), --  9900 / 0x26ac -- last item of row
    1440 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    1441 => std_logic_vector(to_unsigned(  452, 16)), --   452 / 0x01c4
    1442 => std_logic_vector(to_unsigned( 7374, 16)), --  7374 / 0x1cce -- last item of row
    1443 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    1444 => std_logic_vector(to_unsigned(18206, 16)), -- 18206 / 0x471e
    1445 => std_logic_vector(to_unsigned( 9921, 16)), --  9921 / 0x26c1 -- last item of row
    1446 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    1447 => std_logic_vector(to_unsigned( 6131, 16)), --  6131 / 0x17f3
    1448 => std_logic_vector(to_unsigned( 5414, 16)), --  5414 / 0x1526 -- last item of row
    1449 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    1450 => std_logic_vector(to_unsigned(10077, 16)), -- 10077 / 0x275d
    1451 => std_logic_vector(to_unsigned( 9726, 16)), --  9726 / 0x25fe -- last item of row
    1452 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    1453 => std_logic_vector(to_unsigned(12045, 16)), -- 12045 / 0x2f0d
    1454 => std_logic_vector(to_unsigned( 5479, 16)), --  5479 / 0x1567 -- last item of row
    1455 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    1456 => std_logic_vector(to_unsigned( 4322, 16)), --  4322 / 0x10e2
    1457 => std_logic_vector(to_unsigned( 7990, 16)), --  7990 / 0x1f36 -- last item of row
    1458 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    1459 => std_logic_vector(to_unsigned(15616, 16)), -- 15616 / 0x3d00
    1460 => std_logic_vector(to_unsigned( 5550, 16)), --  5550 / 0x15ae -- last item of row
    1461 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    1462 => std_logic_vector(to_unsigned(15561, 16)), -- 15561 / 0x3cc9
    1463 => std_logic_vector(to_unsigned(10661, 16)), -- 10661 / 0x29a5 -- last item of row
    1464 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    1465 => std_logic_vector(to_unsigned(20718, 16)), -- 20718 / 0x50ee
    1466 => std_logic_vector(to_unsigned( 7387, 16)), --  7387 / 0x1cdb -- last item of row
    1467 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    1468 => std_logic_vector(to_unsigned( 2518, 16)), --  2518 / 0x09d6
    1469 => std_logic_vector(to_unsigned(18804, 16)), -- 18804 / 0x4974 -- last item of row
    1470 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    1471 => std_logic_vector(to_unsigned( 8984, 16)), --  8984 / 0x2318
    1472 => std_logic_vector(to_unsigned( 2600, 16)), --  2600 / 0x0a28 -- last item of row
    1473 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    1474 => std_logic_vector(to_unsigned( 6516, 16)), --  6516 / 0x1974
    1475 => std_logic_vector(to_unsigned(17909, 16)), -- 17909 / 0x45f5 -- last item of row
    1476 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    1477 => std_logic_vector(to_unsigned(11148, 16)), -- 11148 / 0x2b8c
    1478 => std_logic_vector(to_unsigned(   98, 16)), --    98 / 0x0062 -- last item of row
    1479 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    1480 => std_logic_vector(to_unsigned(20559, 16)), -- 20559 / 0x504f
    1481 => std_logic_vector(to_unsigned( 3704, 16)), --  3704 / 0x0e78 -- last item of row
    1482 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    1483 => std_logic_vector(to_unsigned( 7510, 16)), --  7510 / 0x1d56
    1484 => std_logic_vector(to_unsigned( 1569, 16)), --  1569 / 0x0621 -- last item of row
    1485 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    1486 => std_logic_vector(to_unsigned(16000, 16)), -- 16000 / 0x3e80
    1487 => std_logic_vector(to_unsigned(11692, 16)), -- 11692 / 0x2dac -- last item of row
    1488 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    1489 => std_logic_vector(to_unsigned( 9147, 16)), --  9147 / 0x23bb
    1490 => std_logic_vector(to_unsigned(10303, 16)), -- 10303 / 0x283f -- last item of row
    1491 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    1492 => std_logic_vector(to_unsigned(16650, 16)), -- 16650 / 0x410a
    1493 => std_logic_vector(to_unsigned(  191, 16)), --   191 / 0x00bf -- last item of row
    1494 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    1495 => std_logic_vector(to_unsigned(15577, 16)), -- 15577 / 0x3cd9
    1496 => std_logic_vector(to_unsigned(18685, 16)), -- 18685 / 0x48fd -- last item of row
    1497 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    1498 => std_logic_vector(to_unsigned(17167, 16)), -- 17167 / 0x430f
    1499 => std_logic_vector(to_unsigned(20917, 16)), -- 20917 / 0x51b5 -- last item of row
    1500 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    1501 => std_logic_vector(to_unsigned( 4256, 16)), --  4256 / 0x10a0
    1502 => std_logic_vector(to_unsigned( 3391, 16)), --  3391 / 0x0d3f -- last item of row
    1503 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    1504 => std_logic_vector(to_unsigned(20092, 16)), -- 20092 / 0x4e7c
    1505 => std_logic_vector(to_unsigned(17219, 16)), -- 17219 / 0x4343 -- last item of row
    1506 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    1507 => std_logic_vector(to_unsigned( 9218, 16)), --  9218 / 0x2402
    1508 => std_logic_vector(to_unsigned( 5056, 16)), --  5056 / 0x13c0 -- last item of row
    1509 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    1510 => std_logic_vector(to_unsigned(18429, 16)), -- 18429 / 0x47fd
    1511 => std_logic_vector(to_unsigned( 8472, 16)), --  8472 / 0x2118 -- last item of row
    1512 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    1513 => std_logic_vector(to_unsigned(12093, 16)), -- 12093 / 0x2f3d
    1514 => std_logic_vector(to_unsigned(20753, 16)), -- 20753 / 0x5111 -- last item of row
    1515 => std_logic_vector(to_unsigned(   45, 16)), --    45 / 0x002d
    1516 => std_logic_vector(to_unsigned(16345, 16)), -- 16345 / 0x3fd9
    1517 => std_logic_vector(to_unsigned(12748, 16)), -- 12748 / 0x31cc -- last item of row
    1518 => std_logic_vector(to_unsigned(   46, 16)), --    46 / 0x002e
    1519 => std_logic_vector(to_unsigned(16023, 16)), -- 16023 / 0x3e97
    1520 => std_logic_vector(to_unsigned(11095, 16)), -- 11095 / 0x2b57 -- last item of row
    1521 => std_logic_vector(to_unsigned(   47, 16)), --    47 / 0x002f
    1522 => std_logic_vector(to_unsigned( 5048, 16)), --  5048 / 0x13b8
    1523 => std_logic_vector(to_unsigned(17595, 16)), -- 17595 / 0x44bb -- last item of row
    1524 => std_logic_vector(to_unsigned(   48, 16)), --    48 / 0x0030
    1525 => std_logic_vector(to_unsigned(18995, 16)), -- 18995 / 0x4a33
    1526 => std_logic_vector(to_unsigned( 4817, 16)), --  4817 / 0x12d1 -- last item of row
    1527 => std_logic_vector(to_unsigned(   49, 16)), --    49 / 0x0031
    1528 => std_logic_vector(to_unsigned(16483, 16)), -- 16483 / 0x4063
    1529 => std_logic_vector(to_unsigned( 3536, 16)), --  3536 / 0x0dd0 -- last item of row
    1530 => std_logic_vector(to_unsigned(   50, 16)), --    50 / 0x0032
    1531 => std_logic_vector(to_unsigned( 1439, 16)), --  1439 / 0x059f
    1532 => std_logic_vector(to_unsigned(16148, 16)), -- 16148 / 0x3f14 -- last item of row
    1533 => std_logic_vector(to_unsigned(   51, 16)), --    51 / 0x0033
    1534 => std_logic_vector(to_unsigned( 3661, 16)), --  3661 / 0x0e4d
    1535 => std_logic_vector(to_unsigned( 3039, 16)), --  3039 / 0x0bdf -- last item of row
    1536 => std_logic_vector(to_unsigned(   52, 16)), --    52 / 0x0034
    1537 => std_logic_vector(to_unsigned(19010, 16)), -- 19010 / 0x4a42
    1538 => std_logic_vector(to_unsigned(18121, 16)), -- 18121 / 0x46c9 -- last item of row
    1539 => std_logic_vector(to_unsigned(   53, 16)), --    53 / 0x0035
    1540 => std_logic_vector(to_unsigned( 8968, 16)), --  8968 / 0x2308
    1541 => std_logic_vector(to_unsigned(11793, 16)), -- 11793 / 0x2e11 -- last item of row
    1542 => std_logic_vector(to_unsigned(   54, 16)), --    54 / 0x0036
    1543 => std_logic_vector(to_unsigned(13427, 16)), -- 13427 / 0x3473
    1544 => std_logic_vector(to_unsigned(18003, 16)), -- 18003 / 0x4653 -- last item of row
    1545 => std_logic_vector(to_unsigned(   55, 16)), --    55 / 0x0037
    1546 => std_logic_vector(to_unsigned( 5303, 16)), --  5303 / 0x14b7
    1547 => std_logic_vector(to_unsigned( 3083, 16)), --  3083 / 0x0c0b -- last item of row
    1548 => std_logic_vector(to_unsigned(   56, 16)), --    56 / 0x0038
    1549 => std_logic_vector(to_unsigned(  531, 16)), --   531 / 0x0213
    1550 => std_logic_vector(to_unsigned(16668, 16)), -- 16668 / 0x411c -- last item of row
    1551 => std_logic_vector(to_unsigned(   57, 16)), --    57 / 0x0039
    1552 => std_logic_vector(to_unsigned( 4771, 16)), --  4771 / 0x12a3
    1553 => std_logic_vector(to_unsigned( 6722, 16)), --  6722 / 0x1a42 -- last item of row
    1554 => std_logic_vector(to_unsigned(   58, 16)), --    58 / 0x003a
    1555 => std_logic_vector(to_unsigned( 5695, 16)), --  5695 / 0x163f
    1556 => std_logic_vector(to_unsigned( 7960, 16)), --  7960 / 0x1f18 -- last item of row
    1557 => std_logic_vector(to_unsigned(   59, 16)), --    59 / 0x003b
    1558 => std_logic_vector(to_unsigned( 3589, 16)), --  3589 / 0x0e05
    1559 => std_logic_vector(to_unsigned(14630, 16)), -- 14630 / 0x3926 -- last item of row
    -- Table for fecframe_normal, C2_5
    1560 => std_logic_vector(to_unsigned(31413, 16)), -- 31413 / 0x7ab5
    1561 => std_logic_vector(to_unsigned(18834, 16)), -- 18834 / 0x4992
    1562 => std_logic_vector(to_unsigned(28884, 16)), -- 28884 / 0x70d4
    1563 => std_logic_vector(to_unsigned(  947, 16)), --   947 / 0x03b3
    1564 => std_logic_vector(to_unsigned(23050, 16)), -- 23050 / 0x5a0a
    1565 => std_logic_vector(to_unsigned(14484, 16)), -- 14484 / 0x3894
    1566 => std_logic_vector(to_unsigned(14809, 16)), -- 14809 / 0x39d9
    1567 => std_logic_vector(to_unsigned( 4968, 16)), --  4968 / 0x1368
    1568 => std_logic_vector(to_unsigned(  455, 16)), --   455 / 0x01c7
    1569 => std_logic_vector(to_unsigned(33659, 16)), -- 33659 / 0x837b
    1570 => std_logic_vector(to_unsigned(16666, 16)), -- 16666 / 0x411a
    1571 => std_logic_vector(to_unsigned(19008, 16)), -- 19008 / 0x4a40 -- last item of row
    1572 => std_logic_vector(to_unsigned(13172, 16)), -- 13172 / 0x3374
    1573 => std_logic_vector(to_unsigned(19939, 16)), -- 19939 / 0x4de3
    1574 => std_logic_vector(to_unsigned(13354, 16)), -- 13354 / 0x342a
    1575 => std_logic_vector(to_unsigned(13719, 16)), -- 13719 / 0x3597
    1576 => std_logic_vector(to_unsigned( 6132, 16)), --  6132 / 0x17f4
    1577 => std_logic_vector(to_unsigned(20086, 16)), -- 20086 / 0x4e76
    1578 => std_logic_vector(to_unsigned(34040, 16)), -- 34040 / 0x84f8
    1579 => std_logic_vector(to_unsigned(13442, 16)), -- 13442 / 0x3482
    1580 => std_logic_vector(to_unsigned(27958, 16)), -- 27958 / 0x6d36
    1581 => std_logic_vector(to_unsigned(16813, 16)), -- 16813 / 0x41ad
    1582 => std_logic_vector(to_unsigned(29619, 16)), -- 29619 / 0x73b3
    1583 => std_logic_vector(to_unsigned(16553, 16)), -- 16553 / 0x40a9 -- last item of row
    1584 => std_logic_vector(to_unsigned( 1499, 16)), --  1499 / 0x05db
    1585 => std_logic_vector(to_unsigned(32075, 16)), -- 32075 / 0x7d4b
    1586 => std_logic_vector(to_unsigned(14962, 16)), -- 14962 / 0x3a72
    1587 => std_logic_vector(to_unsigned(11578, 16)), -- 11578 / 0x2d3a
    1588 => std_logic_vector(to_unsigned(11204, 16)), -- 11204 / 0x2bc4
    1589 => std_logic_vector(to_unsigned( 9217, 16)), --  9217 / 0x2401
    1590 => std_logic_vector(to_unsigned(10485, 16)), -- 10485 / 0x28f5
    1591 => std_logic_vector(to_unsigned(23062, 16)), -- 23062 / 0x5a16
    1592 => std_logic_vector(to_unsigned(30936, 16)), -- 30936 / 0x78d8
    1593 => std_logic_vector(to_unsigned(17892, 16)), -- 17892 / 0x45e4
    1594 => std_logic_vector(to_unsigned(24204, 16)), -- 24204 / 0x5e8c
    1595 => std_logic_vector(to_unsigned(24885, 16)), -- 24885 / 0x6135 -- last item of row
    1596 => std_logic_vector(to_unsigned(32490, 16)), -- 32490 / 0x7eea
    1597 => std_logic_vector(to_unsigned(18086, 16)), -- 18086 / 0x46a6
    1598 => std_logic_vector(to_unsigned(18007, 16)), -- 18007 / 0x4657
    1599 => std_logic_vector(to_unsigned( 4957, 16)), --  4957 / 0x135d
    1600 => std_logic_vector(to_unsigned( 7285, 16)), --  7285 / 0x1c75
    1601 => std_logic_vector(to_unsigned(32073, 16)), -- 32073 / 0x7d49
    1602 => std_logic_vector(to_unsigned(19038, 16)), -- 19038 / 0x4a5e
    1603 => std_logic_vector(to_unsigned( 7152, 16)), --  7152 / 0x1bf0
    1604 => std_logic_vector(to_unsigned(12486, 16)), -- 12486 / 0x30c6
    1605 => std_logic_vector(to_unsigned(13483, 16)), -- 13483 / 0x34ab
    1606 => std_logic_vector(to_unsigned(24808, 16)), -- 24808 / 0x60e8
    1607 => std_logic_vector(to_unsigned(21759, 16)), -- 21759 / 0x54ff -- last item of row
    1608 => std_logic_vector(to_unsigned(32321, 16)), -- 32321 / 0x7e41
    1609 => std_logic_vector(to_unsigned(10839, 16)), -- 10839 / 0x2a57
    1610 => std_logic_vector(to_unsigned(15620, 16)), -- 15620 / 0x3d04
    1611 => std_logic_vector(to_unsigned(33521, 16)), -- 33521 / 0x82f1
    1612 => std_logic_vector(to_unsigned(23030, 16)), -- 23030 / 0x59f6
    1613 => std_logic_vector(to_unsigned(10646, 16)), -- 10646 / 0x2996
    1614 => std_logic_vector(to_unsigned(26236, 16)), -- 26236 / 0x667c
    1615 => std_logic_vector(to_unsigned(19744, 16)), -- 19744 / 0x4d20
    1616 => std_logic_vector(to_unsigned(21713, 16)), -- 21713 / 0x54d1
    1617 => std_logic_vector(to_unsigned(36784, 16)), -- 36784 / 0x8fb0
    1618 => std_logic_vector(to_unsigned( 8016, 16)), --  8016 / 0x1f50
    1619 => std_logic_vector(to_unsigned(12869, 16)), -- 12869 / 0x3245 -- last item of row
    1620 => std_logic_vector(to_unsigned(35597, 16)), -- 35597 / 0x8b0d
    1621 => std_logic_vector(to_unsigned(11129, 16)), -- 11129 / 0x2b79
    1622 => std_logic_vector(to_unsigned(17948, 16)), -- 17948 / 0x461c
    1623 => std_logic_vector(to_unsigned(26160, 16)), -- 26160 / 0x6630
    1624 => std_logic_vector(to_unsigned(14729, 16)), -- 14729 / 0x3989
    1625 => std_logic_vector(to_unsigned(31943, 16)), -- 31943 / 0x7cc7
    1626 => std_logic_vector(to_unsigned(20416, 16)), -- 20416 / 0x4fc0
    1627 => std_logic_vector(to_unsigned(10000, 16)), -- 10000 / 0x2710
    1628 => std_logic_vector(to_unsigned( 7882, 16)), --  7882 / 0x1eca
    1629 => std_logic_vector(to_unsigned(31380, 16)), -- 31380 / 0x7a94
    1630 => std_logic_vector(to_unsigned(27858, 16)), -- 27858 / 0x6cd2
    1631 => std_logic_vector(to_unsigned(33356, 16)), -- 33356 / 0x824c -- last item of row
    1632 => std_logic_vector(to_unsigned(14125, 16)), -- 14125 / 0x372d
    1633 => std_logic_vector(to_unsigned(12131, 16)), -- 12131 / 0x2f63
    1634 => std_logic_vector(to_unsigned(36199, 16)), -- 36199 / 0x8d67
    1635 => std_logic_vector(to_unsigned( 4058, 16)), --  4058 / 0x0fda
    1636 => std_logic_vector(to_unsigned(35992, 16)), -- 35992 / 0x8c98
    1637 => std_logic_vector(to_unsigned(36594, 16)), -- 36594 / 0x8ef2
    1638 => std_logic_vector(to_unsigned(33698, 16)), -- 33698 / 0x83a2
    1639 => std_logic_vector(to_unsigned(15475, 16)), -- 15475 / 0x3c73
    1640 => std_logic_vector(to_unsigned( 1566, 16)), --  1566 / 0x061e
    1641 => std_logic_vector(to_unsigned(18498, 16)), -- 18498 / 0x4842
    1642 => std_logic_vector(to_unsigned(12725, 16)), -- 12725 / 0x31b5
    1643 => std_logic_vector(to_unsigned( 7067, 16)), --  7067 / 0x1b9b -- last item of row
    1644 => std_logic_vector(to_unsigned(17406, 16)), -- 17406 / 0x43fe
    1645 => std_logic_vector(to_unsigned( 8372, 16)), --  8372 / 0x20b4
    1646 => std_logic_vector(to_unsigned(35437, 16)), -- 35437 / 0x8a6d
    1647 => std_logic_vector(to_unsigned( 2888, 16)), --  2888 / 0x0b48
    1648 => std_logic_vector(to_unsigned( 1184, 16)), --  1184 / 0x04a0
    1649 => std_logic_vector(to_unsigned(30068, 16)), -- 30068 / 0x7574
    1650 => std_logic_vector(to_unsigned(25802, 16)), -- 25802 / 0x64ca
    1651 => std_logic_vector(to_unsigned(11056, 16)), -- 11056 / 0x2b30
    1652 => std_logic_vector(to_unsigned( 5507, 16)), --  5507 / 0x1583
    1653 => std_logic_vector(to_unsigned(26313, 16)), -- 26313 / 0x66c9
    1654 => std_logic_vector(to_unsigned(32205, 16)), -- 32205 / 0x7dcd
    1655 => std_logic_vector(to_unsigned(37232, 16)), -- 37232 / 0x9170 -- last item of row
    1656 => std_logic_vector(to_unsigned(15254, 16)), -- 15254 / 0x3b96
    1657 => std_logic_vector(to_unsigned( 5365, 16)), --  5365 / 0x14f5
    1658 => std_logic_vector(to_unsigned(17308, 16)), -- 17308 / 0x439c
    1659 => std_logic_vector(to_unsigned(22519, 16)), -- 22519 / 0x57f7
    1660 => std_logic_vector(to_unsigned(35009, 16)), -- 35009 / 0x88c1
    1661 => std_logic_vector(to_unsigned(  718, 16)), --   718 / 0x02ce
    1662 => std_logic_vector(to_unsigned( 5240, 16)), --  5240 / 0x1478
    1663 => std_logic_vector(to_unsigned(16778, 16)), -- 16778 / 0x418a
    1664 => std_logic_vector(to_unsigned(23131, 16)), -- 23131 / 0x5a5b
    1665 => std_logic_vector(to_unsigned(24092, 16)), -- 24092 / 0x5e1c
    1666 => std_logic_vector(to_unsigned(20587, 16)), -- 20587 / 0x506b
    1667 => std_logic_vector(to_unsigned(33385, 16)), -- 33385 / 0x8269 -- last item of row
    1668 => std_logic_vector(to_unsigned(27455, 16)), -- 27455 / 0x6b3f
    1669 => std_logic_vector(to_unsigned(17602, 16)), -- 17602 / 0x44c2
    1670 => std_logic_vector(to_unsigned( 4590, 16)), --  4590 / 0x11ee
    1671 => std_logic_vector(to_unsigned(21767, 16)), -- 21767 / 0x5507
    1672 => std_logic_vector(to_unsigned(22266, 16)), -- 22266 / 0x56fa
    1673 => std_logic_vector(to_unsigned(27357, 16)), -- 27357 / 0x6add
    1674 => std_logic_vector(to_unsigned(30400, 16)), -- 30400 / 0x76c0
    1675 => std_logic_vector(to_unsigned( 8732, 16)), --  8732 / 0x221c
    1676 => std_logic_vector(to_unsigned( 5596, 16)), --  5596 / 0x15dc
    1677 => std_logic_vector(to_unsigned( 3060, 16)), --  3060 / 0x0bf4
    1678 => std_logic_vector(to_unsigned(33703, 16)), -- 33703 / 0x83a7
    1679 => std_logic_vector(to_unsigned( 3596, 16)), --  3596 / 0x0e0c -- last item of row
    1680 => std_logic_vector(to_unsigned( 6882, 16)), --  6882 / 0x1ae2
    1681 => std_logic_vector(to_unsigned(  873, 16)), --   873 / 0x0369
    1682 => std_logic_vector(to_unsigned(10997, 16)), -- 10997 / 0x2af5
    1683 => std_logic_vector(to_unsigned(24738, 16)), -- 24738 / 0x60a2
    1684 => std_logic_vector(to_unsigned(20770, 16)), -- 20770 / 0x5122
    1685 => std_logic_vector(to_unsigned(10067, 16)), -- 10067 / 0x2753
    1686 => std_logic_vector(to_unsigned(13379, 16)), -- 13379 / 0x3443
    1687 => std_logic_vector(to_unsigned(27409, 16)), -- 27409 / 0x6b11
    1688 => std_logic_vector(to_unsigned(25463, 16)), -- 25463 / 0x6377
    1689 => std_logic_vector(to_unsigned( 2673, 16)), --  2673 / 0x0a71
    1690 => std_logic_vector(to_unsigned( 6998, 16)), --  6998 / 0x1b56
    1691 => std_logic_vector(to_unsigned(31378, 16)), -- 31378 / 0x7a92 -- last item of row
    1692 => std_logic_vector(to_unsigned(15181, 16)), -- 15181 / 0x3b4d
    1693 => std_logic_vector(to_unsigned(13645, 16)), -- 13645 / 0x354d
    1694 => std_logic_vector(to_unsigned(34501, 16)), -- 34501 / 0x86c5
    1695 => std_logic_vector(to_unsigned( 3393, 16)), --  3393 / 0x0d41
    1696 => std_logic_vector(to_unsigned( 3840, 16)), --  3840 / 0x0f00
    1697 => std_logic_vector(to_unsigned(35227, 16)), -- 35227 / 0x899b
    1698 => std_logic_vector(to_unsigned(15562, 16)), -- 15562 / 0x3cca
    1699 => std_logic_vector(to_unsigned(23615, 16)), -- 23615 / 0x5c3f
    1700 => std_logic_vector(to_unsigned(38342, 16)), -- 38342 / 0x95c6
    1701 => std_logic_vector(to_unsigned(12139, 16)), -- 12139 / 0x2f6b
    1702 => std_logic_vector(to_unsigned(19471, 16)), -- 19471 / 0x4c0f
    1703 => std_logic_vector(to_unsigned(15483, 16)), -- 15483 / 0x3c7b -- last item of row
    1704 => std_logic_vector(to_unsigned(13350, 16)), -- 13350 / 0x3426
    1705 => std_logic_vector(to_unsigned( 6707, 16)), --  6707 / 0x1a33
    1706 => std_logic_vector(to_unsigned(23709, 16)), -- 23709 / 0x5c9d
    1707 => std_logic_vector(to_unsigned(37204, 16)), -- 37204 / 0x9154
    1708 => std_logic_vector(to_unsigned(25778, 16)), -- 25778 / 0x64b2
    1709 => std_logic_vector(to_unsigned(21082, 16)), -- 21082 / 0x525a
    1710 => std_logic_vector(to_unsigned( 7511, 16)), --  7511 / 0x1d57
    1711 => std_logic_vector(to_unsigned(14588, 16)), -- 14588 / 0x38fc
    1712 => std_logic_vector(to_unsigned(10010, 16)), -- 10010 / 0x271a
    1713 => std_logic_vector(to_unsigned(21854, 16)), -- 21854 / 0x555e
    1714 => std_logic_vector(to_unsigned(28375, 16)), -- 28375 / 0x6ed7
    1715 => std_logic_vector(to_unsigned(33591, 16)), -- 33591 / 0x8337 -- last item of row
    1716 => std_logic_vector(to_unsigned(12514, 16)), -- 12514 / 0x30e2
    1717 => std_logic_vector(to_unsigned( 4695, 16)), --  4695 / 0x1257
    1718 => std_logic_vector(to_unsigned(37190, 16)), -- 37190 / 0x9146
    1719 => std_logic_vector(to_unsigned(21379, 16)), -- 21379 / 0x5383
    1720 => std_logic_vector(to_unsigned(18723, 16)), -- 18723 / 0x4923
    1721 => std_logic_vector(to_unsigned( 5802, 16)), --  5802 / 0x16aa
    1722 => std_logic_vector(to_unsigned( 7182, 16)), --  7182 / 0x1c0e
    1723 => std_logic_vector(to_unsigned( 2529, 16)), --  2529 / 0x09e1
    1724 => std_logic_vector(to_unsigned(29936, 16)), -- 29936 / 0x74f0
    1725 => std_logic_vector(to_unsigned(35860, 16)), -- 35860 / 0x8c14
    1726 => std_logic_vector(to_unsigned(28338, 16)), -- 28338 / 0x6eb2
    1727 => std_logic_vector(to_unsigned(10835, 16)), -- 10835 / 0x2a53 -- last item of row
    1728 => std_logic_vector(to_unsigned(34283, 16)), -- 34283 / 0x85eb
    1729 => std_logic_vector(to_unsigned(25610, 16)), -- 25610 / 0x640a
    1730 => std_logic_vector(to_unsigned(33026, 16)), -- 33026 / 0x8102
    1731 => std_logic_vector(to_unsigned(31017, 16)), -- 31017 / 0x7929
    1732 => std_logic_vector(to_unsigned(21259, 16)), -- 21259 / 0x530b
    1733 => std_logic_vector(to_unsigned( 2165, 16)), --  2165 / 0x0875
    1734 => std_logic_vector(to_unsigned(21807, 16)), -- 21807 / 0x552f
    1735 => std_logic_vector(to_unsigned(37578, 16)), -- 37578 / 0x92ca
    1736 => std_logic_vector(to_unsigned( 1175, 16)), --  1175 / 0x0497
    1737 => std_logic_vector(to_unsigned(16710, 16)), -- 16710 / 0x4146
    1738 => std_logic_vector(to_unsigned(21939, 16)), -- 21939 / 0x55b3
    1739 => std_logic_vector(to_unsigned(30841, 16)), -- 30841 / 0x7879 -- last item of row
    1740 => std_logic_vector(to_unsigned(27292, 16)), -- 27292 / 0x6a9c
    1741 => std_logic_vector(to_unsigned(33730, 16)), -- 33730 / 0x83c2
    1742 => std_logic_vector(to_unsigned( 6836, 16)), --  6836 / 0x1ab4
    1743 => std_logic_vector(to_unsigned(26476, 16)), -- 26476 / 0x676c
    1744 => std_logic_vector(to_unsigned(27539, 16)), -- 27539 / 0x6b93
    1745 => std_logic_vector(to_unsigned(35784, 16)), -- 35784 / 0x8bc8
    1746 => std_logic_vector(to_unsigned(18245, 16)), -- 18245 / 0x4745
    1747 => std_logic_vector(to_unsigned(16394, 16)), -- 16394 / 0x400a
    1748 => std_logic_vector(to_unsigned(17939, 16)), -- 17939 / 0x4613
    1749 => std_logic_vector(to_unsigned(23094, 16)), -- 23094 / 0x5a36
    1750 => std_logic_vector(to_unsigned(19216, 16)), -- 19216 / 0x4b10
    1751 => std_logic_vector(to_unsigned(17432, 16)), -- 17432 / 0x4418 -- last item of row
    1752 => std_logic_vector(to_unsigned(11655, 16)), -- 11655 / 0x2d87
    1753 => std_logic_vector(to_unsigned( 6183, 16)), --  6183 / 0x1827
    1754 => std_logic_vector(to_unsigned(38708, 16)), -- 38708 / 0x9734
    1755 => std_logic_vector(to_unsigned(28408, 16)), -- 28408 / 0x6ef8
    1756 => std_logic_vector(to_unsigned(35157, 16)), -- 35157 / 0x8955
    1757 => std_logic_vector(to_unsigned(17089, 16)), -- 17089 / 0x42c1
    1758 => std_logic_vector(to_unsigned(13998, 16)), -- 13998 / 0x36ae
    1759 => std_logic_vector(to_unsigned(36029, 16)), -- 36029 / 0x8cbd
    1760 => std_logic_vector(to_unsigned(15052, 16)), -- 15052 / 0x3acc
    1761 => std_logic_vector(to_unsigned(16617, 16)), -- 16617 / 0x40e9
    1762 => std_logic_vector(to_unsigned( 5638, 16)), --  5638 / 0x1606
    1763 => std_logic_vector(to_unsigned(36464, 16)), -- 36464 / 0x8e70 -- last item of row
    1764 => std_logic_vector(to_unsigned(15693, 16)), -- 15693 / 0x3d4d
    1765 => std_logic_vector(to_unsigned(28923, 16)), -- 28923 / 0x70fb
    1766 => std_logic_vector(to_unsigned(26245, 16)), -- 26245 / 0x6685
    1767 => std_logic_vector(to_unsigned( 9432, 16)), --  9432 / 0x24d8
    1768 => std_logic_vector(to_unsigned(11675, 16)), -- 11675 / 0x2d9b
    1769 => std_logic_vector(to_unsigned(25720, 16)), -- 25720 / 0x6478
    1770 => std_logic_vector(to_unsigned(26405, 16)), -- 26405 / 0x6725
    1771 => std_logic_vector(to_unsigned( 5838, 16)), --  5838 / 0x16ce
    1772 => std_logic_vector(to_unsigned(31851, 16)), -- 31851 / 0x7c6b
    1773 => std_logic_vector(to_unsigned(26898, 16)), -- 26898 / 0x6912
    1774 => std_logic_vector(to_unsigned( 8090, 16)), --  8090 / 0x1f9a
    1775 => std_logic_vector(to_unsigned(37037, 16)), -- 37037 / 0x90ad -- last item of row
    1776 => std_logic_vector(to_unsigned(24418, 16)), -- 24418 / 0x5f62
    1777 => std_logic_vector(to_unsigned(27583, 16)), -- 27583 / 0x6bbf
    1778 => std_logic_vector(to_unsigned( 7959, 16)), --  7959 / 0x1f17
    1779 => std_logic_vector(to_unsigned(35562, 16)), -- 35562 / 0x8aea
    1780 => std_logic_vector(to_unsigned(37771, 16)), -- 37771 / 0x938b
    1781 => std_logic_vector(to_unsigned(17784, 16)), -- 17784 / 0x4578
    1782 => std_logic_vector(to_unsigned(11382, 16)), -- 11382 / 0x2c76
    1783 => std_logic_vector(to_unsigned(11156, 16)), -- 11156 / 0x2b94
    1784 => std_logic_vector(to_unsigned(37855, 16)), -- 37855 / 0x93df
    1785 => std_logic_vector(to_unsigned( 7073, 16)), --  7073 / 0x1ba1
    1786 => std_logic_vector(to_unsigned(21685, 16)), -- 21685 / 0x54b5
    1787 => std_logic_vector(to_unsigned(34515, 16)), -- 34515 / 0x86d3 -- last item of row
    1788 => std_logic_vector(to_unsigned(10977, 16)), -- 10977 / 0x2ae1
    1789 => std_logic_vector(to_unsigned(13633, 16)), -- 13633 / 0x3541
    1790 => std_logic_vector(to_unsigned(30969, 16)), -- 30969 / 0x78f9
    1791 => std_logic_vector(to_unsigned( 7516, 16)), --  7516 / 0x1d5c
    1792 => std_logic_vector(to_unsigned(11943, 16)), -- 11943 / 0x2ea7
    1793 => std_logic_vector(to_unsigned(18199, 16)), -- 18199 / 0x4717
    1794 => std_logic_vector(to_unsigned( 5231, 16)), --  5231 / 0x146f
    1795 => std_logic_vector(to_unsigned(13825, 16)), -- 13825 / 0x3601
    1796 => std_logic_vector(to_unsigned(19589, 16)), -- 19589 / 0x4c85
    1797 => std_logic_vector(to_unsigned(23661, 16)), -- 23661 / 0x5c6d
    1798 => std_logic_vector(to_unsigned(11150, 16)), -- 11150 / 0x2b8e
    1799 => std_logic_vector(to_unsigned(35602, 16)), -- 35602 / 0x8b12 -- last item of row
    1800 => std_logic_vector(to_unsigned(19124, 16)), -- 19124 / 0x4ab4
    1801 => std_logic_vector(to_unsigned(30774, 16)), -- 30774 / 0x7836
    1802 => std_logic_vector(to_unsigned( 6670, 16)), --  6670 / 0x1a0e
    1803 => std_logic_vector(to_unsigned(37344, 16)), -- 37344 / 0x91e0
    1804 => std_logic_vector(to_unsigned(16510, 16)), -- 16510 / 0x407e
    1805 => std_logic_vector(to_unsigned(26317, 16)), -- 26317 / 0x66cd
    1806 => std_logic_vector(to_unsigned(23518, 16)), -- 23518 / 0x5bde
    1807 => std_logic_vector(to_unsigned(22957, 16)), -- 22957 / 0x59ad
    1808 => std_logic_vector(to_unsigned( 6348, 16)), --  6348 / 0x18cc
    1809 => std_logic_vector(to_unsigned(34069, 16)), -- 34069 / 0x8515
    1810 => std_logic_vector(to_unsigned( 8845, 16)), --  8845 / 0x228d
    1811 => std_logic_vector(to_unsigned(20175, 16)), -- 20175 / 0x4ecf -- last item of row
    1812 => std_logic_vector(to_unsigned(34985, 16)), -- 34985 / 0x88a9
    1813 => std_logic_vector(to_unsigned(14441, 16)), -- 14441 / 0x3869
    1814 => std_logic_vector(to_unsigned(25668, 16)), -- 25668 / 0x6444
    1815 => std_logic_vector(to_unsigned( 4116, 16)), --  4116 / 0x1014
    1816 => std_logic_vector(to_unsigned( 3019, 16)), --  3019 / 0x0bcb
    1817 => std_logic_vector(to_unsigned(21049, 16)), -- 21049 / 0x5239
    1818 => std_logic_vector(to_unsigned(37308, 16)), -- 37308 / 0x91bc
    1819 => std_logic_vector(to_unsigned(24551, 16)), -- 24551 / 0x5fe7
    1820 => std_logic_vector(to_unsigned(24727, 16)), -- 24727 / 0x6097
    1821 => std_logic_vector(to_unsigned(20104, 16)), -- 20104 / 0x4e88
    1822 => std_logic_vector(to_unsigned(24850, 16)), -- 24850 / 0x6112
    1823 => std_logic_vector(to_unsigned(12114, 16)), -- 12114 / 0x2f52 -- last item of row
    1824 => std_logic_vector(to_unsigned(38187, 16)), -- 38187 / 0x952b
    1825 => std_logic_vector(to_unsigned(28527, 16)), -- 28527 / 0x6f6f
    1826 => std_logic_vector(to_unsigned(13108, 16)), -- 13108 / 0x3334
    1827 => std_logic_vector(to_unsigned(13985, 16)), -- 13985 / 0x36a1
    1828 => std_logic_vector(to_unsigned( 1425, 16)), --  1425 / 0x0591
    1829 => std_logic_vector(to_unsigned(21477, 16)), -- 21477 / 0x53e5
    1830 => std_logic_vector(to_unsigned(30807, 16)), -- 30807 / 0x7857
    1831 => std_logic_vector(to_unsigned( 8613, 16)), --  8613 / 0x21a5
    1832 => std_logic_vector(to_unsigned(26241, 16)), -- 26241 / 0x6681
    1833 => std_logic_vector(to_unsigned(33368, 16)), -- 33368 / 0x8258
    1834 => std_logic_vector(to_unsigned(35913, 16)), -- 35913 / 0x8c49
    1835 => std_logic_vector(to_unsigned(32477, 16)), -- 32477 / 0x7edd -- last item of row
    1836 => std_logic_vector(to_unsigned( 5903, 16)), --  5903 / 0x170f
    1837 => std_logic_vector(to_unsigned(34390, 16)), -- 34390 / 0x8656
    1838 => std_logic_vector(to_unsigned(24641, 16)), -- 24641 / 0x6041
    1839 => std_logic_vector(to_unsigned(26556, 16)), -- 26556 / 0x67bc
    1840 => std_logic_vector(to_unsigned(23007, 16)), -- 23007 / 0x59df
    1841 => std_logic_vector(to_unsigned(27305, 16)), -- 27305 / 0x6aa9
    1842 => std_logic_vector(to_unsigned(38247, 16)), -- 38247 / 0x9567
    1843 => std_logic_vector(to_unsigned( 2621, 16)), --  2621 / 0x0a3d
    1844 => std_logic_vector(to_unsigned( 9122, 16)), --  9122 / 0x23a2
    1845 => std_logic_vector(to_unsigned(32806, 16)), -- 32806 / 0x8026
    1846 => std_logic_vector(to_unsigned(21554, 16)), -- 21554 / 0x5432
    1847 => std_logic_vector(to_unsigned(18685, 16)), -- 18685 / 0x48fd -- last item of row
    1848 => std_logic_vector(to_unsigned(17287, 16)), -- 17287 / 0x4387
    1849 => std_logic_vector(to_unsigned(27292, 16)), -- 27292 / 0x6a9c
    1850 => std_logic_vector(to_unsigned(19033, 16)), -- 19033 / 0x4a59 -- last item of row
    1851 => std_logic_vector(to_unsigned(25796, 16)), -- 25796 / 0x64c4
    1852 => std_logic_vector(to_unsigned(31795, 16)), -- 31795 / 0x7c33
    1853 => std_logic_vector(to_unsigned(12152, 16)), -- 12152 / 0x2f78 -- last item of row
    1854 => std_logic_vector(to_unsigned(12184, 16)), -- 12184 / 0x2f98
    1855 => std_logic_vector(to_unsigned(35088, 16)), -- 35088 / 0x8910
    1856 => std_logic_vector(to_unsigned(31226, 16)), -- 31226 / 0x79fa -- last item of row
    1857 => std_logic_vector(to_unsigned(38263, 16)), -- 38263 / 0x9577
    1858 => std_logic_vector(to_unsigned(33386, 16)), -- 33386 / 0x826a
    1859 => std_logic_vector(to_unsigned(24892, 16)), -- 24892 / 0x613c -- last item of row
    1860 => std_logic_vector(to_unsigned(23114, 16)), -- 23114 / 0x5a4a
    1861 => std_logic_vector(to_unsigned(37995, 16)), -- 37995 / 0x946b
    1862 => std_logic_vector(to_unsigned(29796, 16)), -- 29796 / 0x7464 -- last item of row
    1863 => std_logic_vector(to_unsigned(34336, 16)), -- 34336 / 0x8620
    1864 => std_logic_vector(to_unsigned(10551, 16)), -- 10551 / 0x2937
    1865 => std_logic_vector(to_unsigned(36245, 16)), -- 36245 / 0x8d95 -- last item of row
    1866 => std_logic_vector(to_unsigned(35407, 16)), -- 35407 / 0x8a4f
    1867 => std_logic_vector(to_unsigned(  175, 16)), --   175 / 0x00af
    1868 => std_logic_vector(to_unsigned( 7203, 16)), --  7203 / 0x1c23 -- last item of row
    1869 => std_logic_vector(to_unsigned(14654, 16)), -- 14654 / 0x393e
    1870 => std_logic_vector(to_unsigned(38201, 16)), -- 38201 / 0x9539
    1871 => std_logic_vector(to_unsigned(22605, 16)), -- 22605 / 0x584d -- last item of row
    1872 => std_logic_vector(to_unsigned(28404, 16)), -- 28404 / 0x6ef4
    1873 => std_logic_vector(to_unsigned( 6595, 16)), --  6595 / 0x19c3
    1874 => std_logic_vector(to_unsigned( 1018, 16)), --  1018 / 0x03fa -- last item of row
    1875 => std_logic_vector(to_unsigned(19932, 16)), -- 19932 / 0x4ddc
    1876 => std_logic_vector(to_unsigned( 3524, 16)), --  3524 / 0x0dc4
    1877 => std_logic_vector(to_unsigned(29305, 16)), -- 29305 / 0x7279 -- last item of row
    1878 => std_logic_vector(to_unsigned(31749, 16)), -- 31749 / 0x7c05
    1879 => std_logic_vector(to_unsigned(20247, 16)), -- 20247 / 0x4f17
    1880 => std_logic_vector(to_unsigned( 8128, 16)), --  8128 / 0x1fc0 -- last item of row
    1881 => std_logic_vector(to_unsigned(18026, 16)), -- 18026 / 0x466a
    1882 => std_logic_vector(to_unsigned(36357, 16)), -- 36357 / 0x8e05
    1883 => std_logic_vector(to_unsigned(26735, 16)), -- 26735 / 0x686f -- last item of row
    1884 => std_logic_vector(to_unsigned( 7543, 16)), --  7543 / 0x1d77
    1885 => std_logic_vector(to_unsigned(29767, 16)), -- 29767 / 0x7447
    1886 => std_logic_vector(to_unsigned(13588, 16)), -- 13588 / 0x3514 -- last item of row
    1887 => std_logic_vector(to_unsigned(13333, 16)), -- 13333 / 0x3415
    1888 => std_logic_vector(to_unsigned(25965, 16)), -- 25965 / 0x656d
    1889 => std_logic_vector(to_unsigned( 8463, 16)), --  8463 / 0x210f -- last item of row
    1890 => std_logic_vector(to_unsigned(14504, 16)), -- 14504 / 0x38a8
    1891 => std_logic_vector(to_unsigned(36796, 16)), -- 36796 / 0x8fbc
    1892 => std_logic_vector(to_unsigned(19710, 16)), -- 19710 / 0x4cfe -- last item of row
    1893 => std_logic_vector(to_unsigned( 4528, 16)), --  4528 / 0x11b0
    1894 => std_logic_vector(to_unsigned(25299, 16)), -- 25299 / 0x62d3
    1895 => std_logic_vector(to_unsigned( 7318, 16)), --  7318 / 0x1c96 -- last item of row
    1896 => std_logic_vector(to_unsigned(35091, 16)), -- 35091 / 0x8913
    1897 => std_logic_vector(to_unsigned(25550, 16)), -- 25550 / 0x63ce
    1898 => std_logic_vector(to_unsigned(14798, 16)), -- 14798 / 0x39ce -- last item of row
    1899 => std_logic_vector(to_unsigned( 7824, 16)), --  7824 / 0x1e90
    1900 => std_logic_vector(to_unsigned(  215, 16)), --   215 / 0x00d7
    1901 => std_logic_vector(to_unsigned( 1248, 16)), --  1248 / 0x04e0 -- last item of row
    1902 => std_logic_vector(to_unsigned(30848, 16)), -- 30848 / 0x7880
    1903 => std_logic_vector(to_unsigned( 5362, 16)), --  5362 / 0x14f2
    1904 => std_logic_vector(to_unsigned(17291, 16)), -- 17291 / 0x438b -- last item of row
    1905 => std_logic_vector(to_unsigned(28932, 16)), -- 28932 / 0x7104
    1906 => std_logic_vector(to_unsigned(30249, 16)), -- 30249 / 0x7629
    1907 => std_logic_vector(to_unsigned(27073, 16)), -- 27073 / 0x69c1 -- last item of row
    1908 => std_logic_vector(to_unsigned(13062, 16)), -- 13062 / 0x3306
    1909 => std_logic_vector(to_unsigned( 2103, 16)), --  2103 / 0x0837
    1910 => std_logic_vector(to_unsigned(16206, 16)), -- 16206 / 0x3f4e -- last item of row
    1911 => std_logic_vector(to_unsigned( 7129, 16)), --  7129 / 0x1bd9
    1912 => std_logic_vector(to_unsigned(32062, 16)), -- 32062 / 0x7d3e
    1913 => std_logic_vector(to_unsigned(19612, 16)), -- 19612 / 0x4c9c -- last item of row
    1914 => std_logic_vector(to_unsigned( 9512, 16)), --  9512 / 0x2528
    1915 => std_logic_vector(to_unsigned(21936, 16)), -- 21936 / 0x55b0
    1916 => std_logic_vector(to_unsigned(38833, 16)), -- 38833 / 0x97b1 -- last item of row
    1917 => std_logic_vector(to_unsigned(35849, 16)), -- 35849 / 0x8c09
    1918 => std_logic_vector(to_unsigned(33754, 16)), -- 33754 / 0x83da
    1919 => std_logic_vector(to_unsigned(23450, 16)), -- 23450 / 0x5b9a -- last item of row
    1920 => std_logic_vector(to_unsigned(18705, 16)), -- 18705 / 0x4911
    1921 => std_logic_vector(to_unsigned(28656, 16)), -- 28656 / 0x6ff0
    1922 => std_logic_vector(to_unsigned(18111, 16)), -- 18111 / 0x46bf -- last item of row
    1923 => std_logic_vector(to_unsigned(22749, 16)), -- 22749 / 0x58dd
    1924 => std_logic_vector(to_unsigned(27456, 16)), -- 27456 / 0x6b40
    1925 => std_logic_vector(to_unsigned(32187, 16)), -- 32187 / 0x7dbb -- last item of row
    1926 => std_logic_vector(to_unsigned(28229, 16)), -- 28229 / 0x6e45
    1927 => std_logic_vector(to_unsigned(31684, 16)), -- 31684 / 0x7bc4
    1928 => std_logic_vector(to_unsigned(30160, 16)), -- 30160 / 0x75d0 -- last item of row
    1929 => std_logic_vector(to_unsigned(15293, 16)), -- 15293 / 0x3bbd
    1930 => std_logic_vector(to_unsigned( 8483, 16)), --  8483 / 0x2123
    1931 => std_logic_vector(to_unsigned(28002, 16)), -- 28002 / 0x6d62 -- last item of row
    1932 => std_logic_vector(to_unsigned(14880, 16)), -- 14880 / 0x3a20
    1933 => std_logic_vector(to_unsigned(13334, 16)), -- 13334 / 0x3416
    1934 => std_logic_vector(to_unsigned(12584, 16)), -- 12584 / 0x3128 -- last item of row
    1935 => std_logic_vector(to_unsigned(28646, 16)), -- 28646 / 0x6fe6
    1936 => std_logic_vector(to_unsigned( 2558, 16)), --  2558 / 0x09fe
    1937 => std_logic_vector(to_unsigned(19687, 16)), -- 19687 / 0x4ce7 -- last item of row
    1938 => std_logic_vector(to_unsigned( 6259, 16)), --  6259 / 0x1873
    1939 => std_logic_vector(to_unsigned( 4499, 16)), --  4499 / 0x1193
    1940 => std_logic_vector(to_unsigned(26336, 16)), -- 26336 / 0x66e0 -- last item of row
    1941 => std_logic_vector(to_unsigned(11952, 16)), -- 11952 / 0x2eb0
    1942 => std_logic_vector(to_unsigned(28386, 16)), -- 28386 / 0x6ee2
    1943 => std_logic_vector(to_unsigned( 8405, 16)), --  8405 / 0x20d5 -- last item of row
    1944 => std_logic_vector(to_unsigned(10609, 16)), -- 10609 / 0x2971
    1945 => std_logic_vector(to_unsigned(  961, 16)), --   961 / 0x03c1
    1946 => std_logic_vector(to_unsigned( 7582, 16)), --  7582 / 0x1d9e -- last item of row
    1947 => std_logic_vector(to_unsigned(10423, 16)), -- 10423 / 0x28b7
    1948 => std_logic_vector(to_unsigned(13191, 16)), -- 13191 / 0x3387
    1949 => std_logic_vector(to_unsigned(26818, 16)), -- 26818 / 0x68c2 -- last item of row
    1950 => std_logic_vector(to_unsigned(15922, 16)), -- 15922 / 0x3e32
    1951 => std_logic_vector(to_unsigned(36654, 16)), -- 36654 / 0x8f2e
    1952 => std_logic_vector(to_unsigned(21450, 16)), -- 21450 / 0x53ca -- last item of row
    1953 => std_logic_vector(to_unsigned(10492, 16)), -- 10492 / 0x28fc
    1954 => std_logic_vector(to_unsigned( 1532, 16)), --  1532 / 0x05fc
    1955 => std_logic_vector(to_unsigned( 1205, 16)), --  1205 / 0x04b5 -- last item of row
    1956 => std_logic_vector(to_unsigned(30551, 16)), -- 30551 / 0x7757
    1957 => std_logic_vector(to_unsigned(36482, 16)), -- 36482 / 0x8e82
    1958 => std_logic_vector(to_unsigned(22153, 16)), -- 22153 / 0x5689 -- last item of row
    1959 => std_logic_vector(to_unsigned( 5156, 16)), --  5156 / 0x1424
    1960 => std_logic_vector(to_unsigned(11330, 16)), -- 11330 / 0x2c42
    1961 => std_logic_vector(to_unsigned(34243, 16)), -- 34243 / 0x85c3 -- last item of row
    1962 => std_logic_vector(to_unsigned(28616, 16)), -- 28616 / 0x6fc8
    1963 => std_logic_vector(to_unsigned(35369, 16)), -- 35369 / 0x8a29
    1964 => std_logic_vector(to_unsigned(13322, 16)), -- 13322 / 0x340a -- last item of row
    1965 => std_logic_vector(to_unsigned( 8962, 16)), --  8962 / 0x2302
    1966 => std_logic_vector(to_unsigned( 1485, 16)), --  1485 / 0x05cd
    1967 => std_logic_vector(to_unsigned(21186, 16)), -- 21186 / 0x52c2 -- last item of row
    1968 => std_logic_vector(to_unsigned(23541, 16)), -- 23541 / 0x5bf5
    1969 => std_logic_vector(to_unsigned(17445, 16)), -- 17445 / 0x4425
    1970 => std_logic_vector(to_unsigned(35561, 16)), -- 35561 / 0x8ae9 -- last item of row
    1971 => std_logic_vector(to_unsigned(33133, 16)), -- 33133 / 0x816d
    1972 => std_logic_vector(to_unsigned(11593, 16)), -- 11593 / 0x2d49
    1973 => std_logic_vector(to_unsigned(19895, 16)), -- 19895 / 0x4db7 -- last item of row
    1974 => std_logic_vector(to_unsigned(33917, 16)), -- 33917 / 0x847d
    1975 => std_logic_vector(to_unsigned( 7863, 16)), --  7863 / 0x1eb7
    1976 => std_logic_vector(to_unsigned(33651, 16)), -- 33651 / 0x8373 -- last item of row
    1977 => std_logic_vector(to_unsigned(20063, 16)), -- 20063 / 0x4e5f
    1978 => std_logic_vector(to_unsigned(28331, 16)), -- 28331 / 0x6eab
    1979 => std_logic_vector(to_unsigned(10702, 16)), -- 10702 / 0x29ce -- last item of row
    1980 => std_logic_vector(to_unsigned(13195, 16)), -- 13195 / 0x338b
    1981 => std_logic_vector(to_unsigned(21107, 16)), -- 21107 / 0x5273
    1982 => std_logic_vector(to_unsigned(21859, 16)), -- 21859 / 0x5563 -- last item of row
    1983 => std_logic_vector(to_unsigned( 4364, 16)), --  4364 / 0x110c
    1984 => std_logic_vector(to_unsigned(31137, 16)), -- 31137 / 0x79a1
    1985 => std_logic_vector(to_unsigned( 4804, 16)), --  4804 / 0x12c4 -- last item of row
    1986 => std_logic_vector(to_unsigned( 5585, 16)), --  5585 / 0x15d1
    1987 => std_logic_vector(to_unsigned( 2037, 16)), --  2037 / 0x07f5
    1988 => std_logic_vector(to_unsigned( 4830, 16)), --  4830 / 0x12de -- last item of row
    1989 => std_logic_vector(to_unsigned(30672, 16)), -- 30672 / 0x77d0
    1990 => std_logic_vector(to_unsigned(16927, 16)), -- 16927 / 0x421f
    1991 => std_logic_vector(to_unsigned(14800, 16)), -- 14800 / 0x39d0 -- last item of row
    -- Table for fecframe_normal, C3_4
    1992 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    1993 => std_logic_vector(to_unsigned( 6385, 16)), --  6385 / 0x18f1
    1994 => std_logic_vector(to_unsigned( 7901, 16)), --  7901 / 0x1edd
    1995 => std_logic_vector(to_unsigned(14611, 16)), -- 14611 / 0x3913
    1996 => std_logic_vector(to_unsigned(13389, 16)), -- 13389 / 0x344d
    1997 => std_logic_vector(to_unsigned(11200, 16)), -- 11200 / 0x2bc0
    1998 => std_logic_vector(to_unsigned( 3252, 16)), --  3252 / 0x0cb4
    1999 => std_logic_vector(to_unsigned( 5243, 16)), --  5243 / 0x147b
    2000 => std_logic_vector(to_unsigned( 2504, 16)), --  2504 / 0x09c8
    2001 => std_logic_vector(to_unsigned( 2722, 16)), --  2722 / 0x0aa2
    2002 => std_logic_vector(to_unsigned(  821, 16)), --   821 / 0x0335
    2003 => std_logic_vector(to_unsigned( 7374, 16)), --  7374 / 0x1cce -- last item of row
    2004 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    2005 => std_logic_vector(to_unsigned(11359, 16)), -- 11359 / 0x2c5f
    2006 => std_logic_vector(to_unsigned( 2698, 16)), --  2698 / 0x0a8a
    2007 => std_logic_vector(to_unsigned(  357, 16)), --   357 / 0x0165
    2008 => std_logic_vector(to_unsigned(13824, 16)), -- 13824 / 0x3600
    2009 => std_logic_vector(to_unsigned(12772, 16)), -- 12772 / 0x31e4
    2010 => std_logic_vector(to_unsigned( 7244, 16)), --  7244 / 0x1c4c
    2011 => std_logic_vector(to_unsigned( 6752, 16)), --  6752 / 0x1a60
    2012 => std_logic_vector(to_unsigned(15310, 16)), -- 15310 / 0x3bce
    2013 => std_logic_vector(to_unsigned(  852, 16)), --   852 / 0x0354
    2014 => std_logic_vector(to_unsigned( 2001, 16)), --  2001 / 0x07d1
    2015 => std_logic_vector(to_unsigned(11417, 16)), -- 11417 / 0x2c99 -- last item of row
    2016 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    2017 => std_logic_vector(to_unsigned( 7862, 16)), --  7862 / 0x1eb6
    2018 => std_logic_vector(to_unsigned( 7977, 16)), --  7977 / 0x1f29
    2019 => std_logic_vector(to_unsigned( 6321, 16)), --  6321 / 0x18b1
    2020 => std_logic_vector(to_unsigned(13612, 16)), -- 13612 / 0x352c
    2021 => std_logic_vector(to_unsigned(12197, 16)), -- 12197 / 0x2fa5
    2022 => std_logic_vector(to_unsigned(14449, 16)), -- 14449 / 0x3871
    2023 => std_logic_vector(to_unsigned(15137, 16)), -- 15137 / 0x3b21
    2024 => std_logic_vector(to_unsigned(13860, 16)), -- 13860 / 0x3624
    2025 => std_logic_vector(to_unsigned( 1708, 16)), --  1708 / 0x06ac
    2026 => std_logic_vector(to_unsigned( 6399, 16)), --  6399 / 0x18ff
    2027 => std_logic_vector(to_unsigned(13444, 16)), -- 13444 / 0x3484 -- last item of row
    2028 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    2029 => std_logic_vector(to_unsigned( 1560, 16)), --  1560 / 0x0618
    2030 => std_logic_vector(to_unsigned(11804, 16)), -- 11804 / 0x2e1c
    2031 => std_logic_vector(to_unsigned( 6975, 16)), --  6975 / 0x1b3f
    2032 => std_logic_vector(to_unsigned(13292, 16)), -- 13292 / 0x33ec
    2033 => std_logic_vector(to_unsigned( 3646, 16)), --  3646 / 0x0e3e
    2034 => std_logic_vector(to_unsigned( 3812, 16)), --  3812 / 0x0ee4
    2035 => std_logic_vector(to_unsigned( 8772, 16)), --  8772 / 0x2244
    2036 => std_logic_vector(to_unsigned( 7306, 16)), --  7306 / 0x1c8a
    2037 => std_logic_vector(to_unsigned( 5795, 16)), --  5795 / 0x16a3
    2038 => std_logic_vector(to_unsigned(14327, 16)), -- 14327 / 0x37f7
    2039 => std_logic_vector(to_unsigned( 7866, 16)), --  7866 / 0x1eba -- last item of row
    2040 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    2041 => std_logic_vector(to_unsigned( 7626, 16)), --  7626 / 0x1dca
    2042 => std_logic_vector(to_unsigned(11407, 16)), -- 11407 / 0x2c8f
    2043 => std_logic_vector(to_unsigned(14599, 16)), -- 14599 / 0x3907
    2044 => std_logic_vector(to_unsigned( 9689, 16)), --  9689 / 0x25d9
    2045 => std_logic_vector(to_unsigned( 1628, 16)), --  1628 / 0x065c
    2046 => std_logic_vector(to_unsigned( 2113, 16)), --  2113 / 0x0841
    2047 => std_logic_vector(to_unsigned(10809, 16)), -- 10809 / 0x2a39
    2048 => std_logic_vector(to_unsigned( 9283, 16)), --  9283 / 0x2443
    2049 => std_logic_vector(to_unsigned( 1230, 16)), --  1230 / 0x04ce
    2050 => std_logic_vector(to_unsigned(15241, 16)), -- 15241 / 0x3b89
    2051 => std_logic_vector(to_unsigned( 4870, 16)), --  4870 / 0x1306 -- last item of row
    2052 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    2053 => std_logic_vector(to_unsigned( 1610, 16)), --  1610 / 0x064a
    2054 => std_logic_vector(to_unsigned( 5699, 16)), --  5699 / 0x1643
    2055 => std_logic_vector(to_unsigned(15876, 16)), -- 15876 / 0x3e04
    2056 => std_logic_vector(to_unsigned( 9446, 16)), --  9446 / 0x24e6
    2057 => std_logic_vector(to_unsigned(12515, 16)), -- 12515 / 0x30e3
    2058 => std_logic_vector(to_unsigned( 1400, 16)), --  1400 / 0x0578
    2059 => std_logic_vector(to_unsigned( 6303, 16)), --  6303 / 0x189f
    2060 => std_logic_vector(to_unsigned( 5411, 16)), --  5411 / 0x1523
    2061 => std_logic_vector(to_unsigned(14181, 16)), -- 14181 / 0x3765
    2062 => std_logic_vector(to_unsigned(13925, 16)), -- 13925 / 0x3665
    2063 => std_logic_vector(to_unsigned( 7358, 16)), --  7358 / 0x1cbe -- last item of row
    2064 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    2065 => std_logic_vector(to_unsigned( 4059, 16)), --  4059 / 0x0fdb
    2066 => std_logic_vector(to_unsigned( 8836, 16)), --  8836 / 0x2284
    2067 => std_logic_vector(to_unsigned( 3405, 16)), --  3405 / 0x0d4d
    2068 => std_logic_vector(to_unsigned( 7853, 16)), --  7853 / 0x1ead
    2069 => std_logic_vector(to_unsigned( 7992, 16)), --  7992 / 0x1f38
    2070 => std_logic_vector(to_unsigned(15336, 16)), -- 15336 / 0x3be8
    2071 => std_logic_vector(to_unsigned( 5970, 16)), --  5970 / 0x1752
    2072 => std_logic_vector(to_unsigned(10368, 16)), -- 10368 / 0x2880
    2073 => std_logic_vector(to_unsigned(10278, 16)), -- 10278 / 0x2826
    2074 => std_logic_vector(to_unsigned( 9675, 16)), --  9675 / 0x25cb
    2075 => std_logic_vector(to_unsigned( 4651, 16)), --  4651 / 0x122b -- last item of row
    2076 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    2077 => std_logic_vector(to_unsigned( 4441, 16)), --  4441 / 0x1159
    2078 => std_logic_vector(to_unsigned( 3963, 16)), --  3963 / 0x0f7b
    2079 => std_logic_vector(to_unsigned( 9153, 16)), --  9153 / 0x23c1
    2080 => std_logic_vector(to_unsigned( 2109, 16)), --  2109 / 0x083d
    2081 => std_logic_vector(to_unsigned(12683, 16)), -- 12683 / 0x318b
    2082 => std_logic_vector(to_unsigned( 7459, 16)), --  7459 / 0x1d23
    2083 => std_logic_vector(to_unsigned(12030, 16)), -- 12030 / 0x2efe
    2084 => std_logic_vector(to_unsigned(12221, 16)), -- 12221 / 0x2fbd
    2085 => std_logic_vector(to_unsigned(  629, 16)), --   629 / 0x0275
    2086 => std_logic_vector(to_unsigned(15212, 16)), -- 15212 / 0x3b6c
    2087 => std_logic_vector(to_unsigned(  406, 16)), --   406 / 0x0196 -- last item of row
    2088 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    2089 => std_logic_vector(to_unsigned( 6007, 16)), --  6007 / 0x1777
    2090 => std_logic_vector(to_unsigned( 8411, 16)), --  8411 / 0x20db
    2091 => std_logic_vector(to_unsigned( 5771, 16)), --  5771 / 0x168b
    2092 => std_logic_vector(to_unsigned( 3497, 16)), --  3497 / 0x0da9
    2093 => std_logic_vector(to_unsigned(  543, 16)), --   543 / 0x021f
    2094 => std_logic_vector(to_unsigned(14202, 16)), -- 14202 / 0x377a
    2095 => std_logic_vector(to_unsigned(  875, 16)), --   875 / 0x036b
    2096 => std_logic_vector(to_unsigned( 9186, 16)), --  9186 / 0x23e2
    2097 => std_logic_vector(to_unsigned( 6235, 16)), --  6235 / 0x185b
    2098 => std_logic_vector(to_unsigned(13908, 16)), -- 13908 / 0x3654
    2099 => std_logic_vector(to_unsigned( 3563, 16)), --  3563 / 0x0deb -- last item of row
    2100 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    2101 => std_logic_vector(to_unsigned( 3232, 16)), --  3232 / 0x0ca0
    2102 => std_logic_vector(to_unsigned( 6625, 16)), --  6625 / 0x19e1
    2103 => std_logic_vector(to_unsigned( 4795, 16)), --  4795 / 0x12bb
    2104 => std_logic_vector(to_unsigned(  546, 16)), --   546 / 0x0222
    2105 => std_logic_vector(to_unsigned( 9781, 16)), --  9781 / 0x2635
    2106 => std_logic_vector(to_unsigned( 2071, 16)), --  2071 / 0x0817
    2107 => std_logic_vector(to_unsigned( 7312, 16)), --  7312 / 0x1c90
    2108 => std_logic_vector(to_unsigned( 3399, 16)), --  3399 / 0x0d47
    2109 => std_logic_vector(to_unsigned( 7250, 16)), --  7250 / 0x1c52
    2110 => std_logic_vector(to_unsigned( 4932, 16)), --  4932 / 0x1344
    2111 => std_logic_vector(to_unsigned(12652, 16)), -- 12652 / 0x316c -- last item of row
    2112 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    2113 => std_logic_vector(to_unsigned( 8820, 16)), --  8820 / 0x2274
    2114 => std_logic_vector(to_unsigned(10088, 16)), -- 10088 / 0x2768
    2115 => std_logic_vector(to_unsigned(11090, 16)), -- 11090 / 0x2b52
    2116 => std_logic_vector(to_unsigned( 7069, 16)), --  7069 / 0x1b9d
    2117 => std_logic_vector(to_unsigned( 6585, 16)), --  6585 / 0x19b9
    2118 => std_logic_vector(to_unsigned(13134, 16)), -- 13134 / 0x334e
    2119 => std_logic_vector(to_unsigned(10158, 16)), -- 10158 / 0x27ae
    2120 => std_logic_vector(to_unsigned( 7183, 16)), --  7183 / 0x1c0f
    2121 => std_logic_vector(to_unsigned(  488, 16)), --   488 / 0x01e8
    2122 => std_logic_vector(to_unsigned( 7455, 16)), --  7455 / 0x1d1f
    2123 => std_logic_vector(to_unsigned( 9238, 16)), --  9238 / 0x2416 -- last item of row
    2124 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    2125 => std_logic_vector(to_unsigned( 1903, 16)), --  1903 / 0x076f
    2126 => std_logic_vector(to_unsigned(10818, 16)), -- 10818 / 0x2a42
    2127 => std_logic_vector(to_unsigned(  119, 16)), --   119 / 0x0077
    2128 => std_logic_vector(to_unsigned(  215, 16)), --   215 / 0x00d7
    2129 => std_logic_vector(to_unsigned( 7558, 16)), --  7558 / 0x1d86
    2130 => std_logic_vector(to_unsigned(11046, 16)), -- 11046 / 0x2b26
    2131 => std_logic_vector(to_unsigned(10615, 16)), -- 10615 / 0x2977
    2132 => std_logic_vector(to_unsigned(11545, 16)), -- 11545 / 0x2d19
    2133 => std_logic_vector(to_unsigned(14784, 16)), -- 14784 / 0x39c0
    2134 => std_logic_vector(to_unsigned( 7961, 16)), --  7961 / 0x1f19
    2135 => std_logic_vector(to_unsigned(15619, 16)), -- 15619 / 0x3d03 -- last item of row
    2136 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    2137 => std_logic_vector(to_unsigned( 3655, 16)), --  3655 / 0x0e47
    2138 => std_logic_vector(to_unsigned( 8736, 16)), --  8736 / 0x2220
    2139 => std_logic_vector(to_unsigned( 4917, 16)), --  4917 / 0x1335
    2140 => std_logic_vector(to_unsigned(15874, 16)), -- 15874 / 0x3e02
    2141 => std_logic_vector(to_unsigned( 5129, 16)), --  5129 / 0x1409
    2142 => std_logic_vector(to_unsigned( 2134, 16)), --  2134 / 0x0856
    2143 => std_logic_vector(to_unsigned(15944, 16)), -- 15944 / 0x3e48
    2144 => std_logic_vector(to_unsigned(14768, 16)), -- 14768 / 0x39b0
    2145 => std_logic_vector(to_unsigned( 7150, 16)), --  7150 / 0x1bee
    2146 => std_logic_vector(to_unsigned( 2692, 16)), --  2692 / 0x0a84
    2147 => std_logic_vector(to_unsigned( 1469, 16)), --  1469 / 0x05bd -- last item of row
    2148 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    2149 => std_logic_vector(to_unsigned( 8316, 16)), --  8316 / 0x207c
    2150 => std_logic_vector(to_unsigned( 3820, 16)), --  3820 / 0x0eec
    2151 => std_logic_vector(to_unsigned(  505, 16)), --   505 / 0x01f9
    2152 => std_logic_vector(to_unsigned( 8923, 16)), --  8923 / 0x22db
    2153 => std_logic_vector(to_unsigned( 6757, 16)), --  6757 / 0x1a65
    2154 => std_logic_vector(to_unsigned(  806, 16)), --   806 / 0x0326
    2155 => std_logic_vector(to_unsigned( 7957, 16)), --  7957 / 0x1f15
    2156 => std_logic_vector(to_unsigned( 4216, 16)), --  4216 / 0x1078
    2157 => std_logic_vector(to_unsigned(15589, 16)), -- 15589 / 0x3ce5
    2158 => std_logic_vector(to_unsigned(13244, 16)), -- 13244 / 0x33bc
    2159 => std_logic_vector(to_unsigned( 2622, 16)), --  2622 / 0x0a3e -- last item of row
    2160 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    2161 => std_logic_vector(to_unsigned(14463, 16)), -- 14463 / 0x387f
    2162 => std_logic_vector(to_unsigned( 4852, 16)), --  4852 / 0x12f4
    2163 => std_logic_vector(to_unsigned(15733, 16)), -- 15733 / 0x3d75
    2164 => std_logic_vector(to_unsigned( 3041, 16)), --  3041 / 0x0be1
    2165 => std_logic_vector(to_unsigned(11193, 16)), -- 11193 / 0x2bb9
    2166 => std_logic_vector(to_unsigned(12860, 16)), -- 12860 / 0x323c
    2167 => std_logic_vector(to_unsigned(13673, 16)), -- 13673 / 0x3569
    2168 => std_logic_vector(to_unsigned( 8152, 16)), --  8152 / 0x1fd8
    2169 => std_logic_vector(to_unsigned( 6551, 16)), --  6551 / 0x1997
    2170 => std_logic_vector(to_unsigned(15108, 16)), -- 15108 / 0x3b04
    2171 => std_logic_vector(to_unsigned( 8758, 16)), --  8758 / 0x2236 -- last item of row
    2172 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    2173 => std_logic_vector(to_unsigned( 3149, 16)), --  3149 / 0x0c4d
    2174 => std_logic_vector(to_unsigned(11981, 16)), -- 11981 / 0x2ecd -- last item of row
    2175 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    2176 => std_logic_vector(to_unsigned(13416, 16)), -- 13416 / 0x3468
    2177 => std_logic_vector(to_unsigned( 6906, 16)), --  6906 / 0x1afa -- last item of row
    2178 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    2179 => std_logic_vector(to_unsigned(13098, 16)), -- 13098 / 0x332a
    2180 => std_logic_vector(to_unsigned(13352, 16)), -- 13352 / 0x3428 -- last item of row
    2181 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    2182 => std_logic_vector(to_unsigned( 2009, 16)), --  2009 / 0x07d9
    2183 => std_logic_vector(to_unsigned(14460, 16)), -- 14460 / 0x387c -- last item of row
    2184 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    2185 => std_logic_vector(to_unsigned( 7207, 16)), --  7207 / 0x1c27
    2186 => std_logic_vector(to_unsigned( 4314, 16)), --  4314 / 0x10da -- last item of row
    2187 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    2188 => std_logic_vector(to_unsigned( 3312, 16)), --  3312 / 0x0cf0
    2189 => std_logic_vector(to_unsigned( 3945, 16)), --  3945 / 0x0f69 -- last item of row
    2190 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    2191 => std_logic_vector(to_unsigned( 4418, 16)), --  4418 / 0x1142
    2192 => std_logic_vector(to_unsigned( 6248, 16)), --  6248 / 0x1868 -- last item of row
    2193 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    2194 => std_logic_vector(to_unsigned( 2669, 16)), --  2669 / 0x0a6d
    2195 => std_logic_vector(to_unsigned(13975, 16)), -- 13975 / 0x3697 -- last item of row
    2196 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    2197 => std_logic_vector(to_unsigned( 7571, 16)), --  7571 / 0x1d93
    2198 => std_logic_vector(to_unsigned( 9023, 16)), --  9023 / 0x233f -- last item of row
    2199 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    2200 => std_logic_vector(to_unsigned(14172, 16)), -- 14172 / 0x375c
    2201 => std_logic_vector(to_unsigned( 2967, 16)), --  2967 / 0x0b97 -- last item of row
    2202 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    2203 => std_logic_vector(to_unsigned( 7271, 16)), --  7271 / 0x1c67
    2204 => std_logic_vector(to_unsigned( 7138, 16)), --  7138 / 0x1be2 -- last item of row
    2205 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    2206 => std_logic_vector(to_unsigned( 6135, 16)), --  6135 / 0x17f7
    2207 => std_logic_vector(to_unsigned(13670, 16)), -- 13670 / 0x3566 -- last item of row
    2208 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    2209 => std_logic_vector(to_unsigned( 7490, 16)), --  7490 / 0x1d42
    2210 => std_logic_vector(to_unsigned(14559, 16)), -- 14559 / 0x38df -- last item of row
    2211 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    2212 => std_logic_vector(to_unsigned( 8657, 16)), --  8657 / 0x21d1
    2213 => std_logic_vector(to_unsigned( 2466, 16)), --  2466 / 0x09a2 -- last item of row
    2214 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    2215 => std_logic_vector(to_unsigned( 8599, 16)), --  8599 / 0x2197
    2216 => std_logic_vector(to_unsigned(12834, 16)), -- 12834 / 0x3222 -- last item of row
    2217 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    2218 => std_logic_vector(to_unsigned( 3470, 16)), --  3470 / 0x0d8e
    2219 => std_logic_vector(to_unsigned( 3152, 16)), --  3152 / 0x0c50 -- last item of row
    2220 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    2221 => std_logic_vector(to_unsigned(13917, 16)), -- 13917 / 0x365d
    2222 => std_logic_vector(to_unsigned( 4365, 16)), --  4365 / 0x110d -- last item of row
    2223 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    2224 => std_logic_vector(to_unsigned( 6024, 16)), --  6024 / 0x1788
    2225 => std_logic_vector(to_unsigned(13730, 16)), -- 13730 / 0x35a2 -- last item of row
    2226 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    2227 => std_logic_vector(to_unsigned(10973, 16)), -- 10973 / 0x2add
    2228 => std_logic_vector(to_unsigned(14182, 16)), -- 14182 / 0x3766 -- last item of row
    2229 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    2230 => std_logic_vector(to_unsigned( 2464, 16)), --  2464 / 0x09a0
    2231 => std_logic_vector(to_unsigned(13167, 16)), -- 13167 / 0x336f -- last item of row
    2232 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    2233 => std_logic_vector(to_unsigned( 5281, 16)), --  5281 / 0x14a1
    2234 => std_logic_vector(to_unsigned(15049, 16)), -- 15049 / 0x3ac9 -- last item of row
    2235 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    2236 => std_logic_vector(to_unsigned( 1103, 16)), --  1103 / 0x044f
    2237 => std_logic_vector(to_unsigned( 1849, 16)), --  1849 / 0x0739 -- last item of row
    2238 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    2239 => std_logic_vector(to_unsigned( 2058, 16)), --  2058 / 0x080a
    2240 => std_logic_vector(to_unsigned( 1069, 16)), --  1069 / 0x042d -- last item of row
    2241 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    2242 => std_logic_vector(to_unsigned( 9654, 16)), --  9654 / 0x25b6
    2243 => std_logic_vector(to_unsigned( 6095, 16)), --  6095 / 0x17cf -- last item of row
    2244 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    2245 => std_logic_vector(to_unsigned(14311, 16)), -- 14311 / 0x37e7
    2246 => std_logic_vector(to_unsigned( 7667, 16)), --  7667 / 0x1df3 -- last item of row
    2247 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    2248 => std_logic_vector(to_unsigned(15617, 16)), -- 15617 / 0x3d01
    2249 => std_logic_vector(to_unsigned( 8146, 16)), --  8146 / 0x1fd2 -- last item of row
    2250 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    2251 => std_logic_vector(to_unsigned( 4588, 16)), --  4588 / 0x11ec
    2252 => std_logic_vector(to_unsigned(11218, 16)), -- 11218 / 0x2bd2 -- last item of row
    2253 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    2254 => std_logic_vector(to_unsigned(13660, 16)), -- 13660 / 0x355c
    2255 => std_logic_vector(to_unsigned( 6243, 16)), --  6243 / 0x1863 -- last item of row
    2256 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    2257 => std_logic_vector(to_unsigned( 8578, 16)), --  8578 / 0x2182
    2258 => std_logic_vector(to_unsigned( 7874, 16)), --  7874 / 0x1ec2 -- last item of row
    2259 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    2260 => std_logic_vector(to_unsigned(11741, 16)), -- 11741 / 0x2ddd
    2261 => std_logic_vector(to_unsigned( 2686, 16)), --  2686 / 0x0a7e -- last item of row
    2262 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    2263 => std_logic_vector(to_unsigned( 1022, 16)), --  1022 / 0x03fe
    2264 => std_logic_vector(to_unsigned( 1264, 16)), --  1264 / 0x04f0 -- last item of row
    2265 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    2266 => std_logic_vector(to_unsigned(12604, 16)), -- 12604 / 0x313c
    2267 => std_logic_vector(to_unsigned( 9965, 16)), --  9965 / 0x26ed -- last item of row
    2268 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    2269 => std_logic_vector(to_unsigned( 8217, 16)), --  8217 / 0x2019
    2270 => std_logic_vector(to_unsigned( 2707, 16)), --  2707 / 0x0a93 -- last item of row
    2271 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    2272 => std_logic_vector(to_unsigned( 3156, 16)), --  3156 / 0x0c54
    2273 => std_logic_vector(to_unsigned(11793, 16)), -- 11793 / 0x2e11 -- last item of row
    2274 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    2275 => std_logic_vector(to_unsigned(  354, 16)), --   354 / 0x0162
    2276 => std_logic_vector(to_unsigned( 1514, 16)), --  1514 / 0x05ea -- last item of row
    2277 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    2278 => std_logic_vector(to_unsigned( 6978, 16)), --  6978 / 0x1b42
    2279 => std_logic_vector(to_unsigned(14058, 16)), -- 14058 / 0x36ea -- last item of row
    2280 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    2281 => std_logic_vector(to_unsigned( 7922, 16)), --  7922 / 0x1ef2
    2282 => std_logic_vector(to_unsigned(16079, 16)), -- 16079 / 0x3ecf -- last item of row
    2283 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    2284 => std_logic_vector(to_unsigned(15087, 16)), -- 15087 / 0x3aef
    2285 => std_logic_vector(to_unsigned(12138, 16)), -- 12138 / 0x2f6a -- last item of row
    2286 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    2287 => std_logic_vector(to_unsigned( 5053, 16)), --  5053 / 0x13bd
    2288 => std_logic_vector(to_unsigned( 6470, 16)), --  6470 / 0x1946 -- last item of row
    2289 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    2290 => std_logic_vector(to_unsigned(12687, 16)), -- 12687 / 0x318f
    2291 => std_logic_vector(to_unsigned(14932, 16)), -- 14932 / 0x3a54 -- last item of row
    2292 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    2293 => std_logic_vector(to_unsigned(15458, 16)), -- 15458 / 0x3c62
    2294 => std_logic_vector(to_unsigned( 1763, 16)), --  1763 / 0x06e3 -- last item of row
    2295 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    2296 => std_logic_vector(to_unsigned( 8121, 16)), --  8121 / 0x1fb9
    2297 => std_logic_vector(to_unsigned( 1721, 16)), --  1721 / 0x06b9 -- last item of row
    2298 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    2299 => std_logic_vector(to_unsigned(12431, 16)), -- 12431 / 0x308f
    2300 => std_logic_vector(to_unsigned(  549, 16)), --   549 / 0x0225 -- last item of row
    2301 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    2302 => std_logic_vector(to_unsigned( 4129, 16)), --  4129 / 0x1021
    2303 => std_logic_vector(to_unsigned( 7091, 16)), --  7091 / 0x1bb3 -- last item of row
    2304 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    2305 => std_logic_vector(to_unsigned( 1426, 16)), --  1426 / 0x0592
    2306 => std_logic_vector(to_unsigned( 8415, 16)), --  8415 / 0x20df -- last item of row
    2307 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    2308 => std_logic_vector(to_unsigned( 9783, 16)), --  9783 / 0x2637
    2309 => std_logic_vector(to_unsigned( 7604, 16)), --  7604 / 0x1db4 -- last item of row
    2310 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    2311 => std_logic_vector(to_unsigned( 6295, 16)), --  6295 / 0x1897
    2312 => std_logic_vector(to_unsigned(11329, 16)), -- 11329 / 0x2c41 -- last item of row
    2313 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    2314 => std_logic_vector(to_unsigned( 1409, 16)), --  1409 / 0x0581
    2315 => std_logic_vector(to_unsigned(12061, 16)), -- 12061 / 0x2f1d -- last item of row
    2316 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    2317 => std_logic_vector(to_unsigned( 8065, 16)), --  8065 / 0x1f81
    2318 => std_logic_vector(to_unsigned( 9087, 16)), --  9087 / 0x237f -- last item of row
    2319 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    2320 => std_logic_vector(to_unsigned( 2918, 16)), --  2918 / 0x0b66
    2321 => std_logic_vector(to_unsigned( 8438, 16)), --  8438 / 0x20f6 -- last item of row
    2322 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    2323 => std_logic_vector(to_unsigned( 1293, 16)), --  1293 / 0x050d
    2324 => std_logic_vector(to_unsigned(14115, 16)), -- 14115 / 0x3723 -- last item of row
    2325 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    2326 => std_logic_vector(to_unsigned( 3922, 16)), --  3922 / 0x0f52
    2327 => std_logic_vector(to_unsigned(13851, 16)), -- 13851 / 0x361b -- last item of row
    2328 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    2329 => std_logic_vector(to_unsigned( 3851, 16)), --  3851 / 0x0f0b
    2330 => std_logic_vector(to_unsigned( 4000, 16)), --  4000 / 0x0fa0 -- last item of row
    2331 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    2332 => std_logic_vector(to_unsigned( 5865, 16)), --  5865 / 0x16e9
    2333 => std_logic_vector(to_unsigned( 1768, 16)), --  1768 / 0x06e8 -- last item of row
    2334 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    2335 => std_logic_vector(to_unsigned( 2655, 16)), --  2655 / 0x0a5f
    2336 => std_logic_vector(to_unsigned(14957, 16)), -- 14957 / 0x3a6d -- last item of row
    2337 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    2338 => std_logic_vector(to_unsigned( 5565, 16)), --  5565 / 0x15bd
    2339 => std_logic_vector(to_unsigned( 6332, 16)), --  6332 / 0x18bc -- last item of row
    2340 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    2341 => std_logic_vector(to_unsigned( 4303, 16)), --  4303 / 0x10cf
    2342 => std_logic_vector(to_unsigned(12631, 16)), -- 12631 / 0x3157 -- last item of row
    2343 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    2344 => std_logic_vector(to_unsigned(11653, 16)), -- 11653 / 0x2d85
    2345 => std_logic_vector(to_unsigned(12236, 16)), -- 12236 / 0x2fcc -- last item of row
    2346 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    2347 => std_logic_vector(to_unsigned(16025, 16)), -- 16025 / 0x3e99
    2348 => std_logic_vector(to_unsigned( 7632, 16)), --  7632 / 0x1dd0 -- last item of row
    2349 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    2350 => std_logic_vector(to_unsigned( 4655, 16)), --  4655 / 0x122f
    2351 => std_logic_vector(to_unsigned(14128, 16)), -- 14128 / 0x3730 -- last item of row
    2352 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    2353 => std_logic_vector(to_unsigned( 9584, 16)), --  9584 / 0x2570
    2354 => std_logic_vector(to_unsigned(13123, 16)), -- 13123 / 0x3343 -- last item of row
    2355 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    2356 => std_logic_vector(to_unsigned(13987, 16)), -- 13987 / 0x36a3
    2357 => std_logic_vector(to_unsigned( 9597, 16)), --  9597 / 0x257d -- last item of row
    2358 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    2359 => std_logic_vector(to_unsigned(15409, 16)), -- 15409 / 0x3c31
    2360 => std_logic_vector(to_unsigned(12110, 16)), -- 12110 / 0x2f4e -- last item of row
    2361 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    2362 => std_logic_vector(to_unsigned( 8754, 16)), --  8754 / 0x2232
    2363 => std_logic_vector(to_unsigned(15490, 16)), -- 15490 / 0x3c82 -- last item of row
    2364 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    2365 => std_logic_vector(to_unsigned( 7416, 16)), --  7416 / 0x1cf8
    2366 => std_logic_vector(to_unsigned(15325, 16)), -- 15325 / 0x3bdd -- last item of row
    2367 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    2368 => std_logic_vector(to_unsigned( 2909, 16)), --  2909 / 0x0b5d
    2369 => std_logic_vector(to_unsigned(15549, 16)), -- 15549 / 0x3cbd -- last item of row
    2370 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    2371 => std_logic_vector(to_unsigned( 2995, 16)), --  2995 / 0x0bb3
    2372 => std_logic_vector(to_unsigned( 8257, 16)), --  8257 / 0x2041 -- last item of row
    2373 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    2374 => std_logic_vector(to_unsigned( 9406, 16)), --  9406 / 0x24be
    2375 => std_logic_vector(to_unsigned( 4791, 16)), --  4791 / 0x12b7 -- last item of row
    2376 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    2377 => std_logic_vector(to_unsigned(11111, 16)), -- 11111 / 0x2b67
    2378 => std_logic_vector(to_unsigned( 4854, 16)), --  4854 / 0x12f6 -- last item of row
    2379 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    2380 => std_logic_vector(to_unsigned( 2812, 16)), --  2812 / 0x0afc
    2381 => std_logic_vector(to_unsigned( 8521, 16)), --  8521 / 0x2149 -- last item of row
    2382 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    2383 => std_logic_vector(to_unsigned( 8476, 16)), --  8476 / 0x211c
    2384 => std_logic_vector(to_unsigned(14717, 16)), -- 14717 / 0x397d -- last item of row
    2385 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    2386 => std_logic_vector(to_unsigned( 7820, 16)), --  7820 / 0x1e8c
    2387 => std_logic_vector(to_unsigned(15360, 16)), -- 15360 / 0x3c00 -- last item of row
    2388 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    2389 => std_logic_vector(to_unsigned( 1179, 16)), --  1179 / 0x049b
    2390 => std_logic_vector(to_unsigned( 7939, 16)), --  7939 / 0x1f03 -- last item of row
    2391 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    2392 => std_logic_vector(to_unsigned( 2357, 16)), --  2357 / 0x0935
    2393 => std_logic_vector(to_unsigned( 8678, 16)), --  8678 / 0x21e6 -- last item of row
    2394 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    2395 => std_logic_vector(to_unsigned( 7703, 16)), --  7703 / 0x1e17
    2396 => std_logic_vector(to_unsigned( 6216, 16)), --  6216 / 0x1848 -- last item of row
    2397 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    2398 => std_logic_vector(to_unsigned( 3477, 16)), --  3477 / 0x0d95
    2399 => std_logic_vector(to_unsigned( 7067, 16)), --  7067 / 0x1b9b -- last item of row
    2400 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    2401 => std_logic_vector(to_unsigned( 3931, 16)), --  3931 / 0x0f5b
    2402 => std_logic_vector(to_unsigned(13845, 16)), -- 13845 / 0x3615 -- last item of row
    2403 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    2404 => std_logic_vector(to_unsigned( 7675, 16)), --  7675 / 0x1dfb
    2405 => std_logic_vector(to_unsigned(12899, 16)), -- 12899 / 0x3263 -- last item of row
    2406 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    2407 => std_logic_vector(to_unsigned( 1754, 16)), --  1754 / 0x06da
    2408 => std_logic_vector(to_unsigned( 8187, 16)), --  8187 / 0x1ffb -- last item of row
    2409 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    2410 => std_logic_vector(to_unsigned( 7785, 16)), --  7785 / 0x1e69
    2411 => std_logic_vector(to_unsigned( 1400, 16)), --  1400 / 0x0578 -- last item of row
    2412 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    2413 => std_logic_vector(to_unsigned( 9213, 16)), --  9213 / 0x23fd
    2414 => std_logic_vector(to_unsigned( 5891, 16)), --  5891 / 0x1703 -- last item of row
    2415 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    2416 => std_logic_vector(to_unsigned( 2494, 16)), --  2494 / 0x09be
    2417 => std_logic_vector(to_unsigned( 7703, 16)), --  7703 / 0x1e17 -- last item of row
    2418 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    2419 => std_logic_vector(to_unsigned( 2576, 16)), --  2576 / 0x0a10
    2420 => std_logic_vector(to_unsigned( 7902, 16)), --  7902 / 0x1ede -- last item of row
    2421 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    2422 => std_logic_vector(to_unsigned( 4821, 16)), --  4821 / 0x12d5
    2423 => std_logic_vector(to_unsigned(15682, 16)), -- 15682 / 0x3d42 -- last item of row
    2424 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    2425 => std_logic_vector(to_unsigned(10426, 16)), -- 10426 / 0x28ba
    2426 => std_logic_vector(to_unsigned(11935, 16)), -- 11935 / 0x2e9f -- last item of row
    2427 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    2428 => std_logic_vector(to_unsigned( 1810, 16)), --  1810 / 0x0712
    2429 => std_logic_vector(to_unsigned(  904, 16)), --   904 / 0x0388 -- last item of row
    2430 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    2431 => std_logic_vector(to_unsigned(11332, 16)), -- 11332 / 0x2c44
    2432 => std_logic_vector(to_unsigned( 9264, 16)), --  9264 / 0x2430 -- last item of row
    2433 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    2434 => std_logic_vector(to_unsigned(11312, 16)), -- 11312 / 0x2c30
    2435 => std_logic_vector(to_unsigned( 3570, 16)), --  3570 / 0x0df2 -- last item of row
    2436 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    2437 => std_logic_vector(to_unsigned(14916, 16)), -- 14916 / 0x3a44
    2438 => std_logic_vector(to_unsigned( 2650, 16)), --  2650 / 0x0a5a -- last item of row
    2439 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    2440 => std_logic_vector(to_unsigned( 7679, 16)), --  7679 / 0x1dff
    2441 => std_logic_vector(to_unsigned( 7842, 16)), --  7842 / 0x1ea2 -- last item of row
    2442 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    2443 => std_logic_vector(to_unsigned( 6089, 16)), --  6089 / 0x17c9
    2444 => std_logic_vector(to_unsigned(13084, 16)), -- 13084 / 0x331c -- last item of row
    2445 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    2446 => std_logic_vector(to_unsigned( 3938, 16)), --  3938 / 0x0f62
    2447 => std_logic_vector(to_unsigned( 2751, 16)), --  2751 / 0x0abf -- last item of row
    2448 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    2449 => std_logic_vector(to_unsigned( 8509, 16)), --  8509 / 0x213d
    2450 => std_logic_vector(to_unsigned( 4648, 16)), --  4648 / 0x1228 -- last item of row
    2451 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    2452 => std_logic_vector(to_unsigned(12204, 16)), -- 12204 / 0x2fac
    2453 => std_logic_vector(to_unsigned( 8917, 16)), --  8917 / 0x22d5 -- last item of row
    2454 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    2455 => std_logic_vector(to_unsigned( 5749, 16)), --  5749 / 0x1675
    2456 => std_logic_vector(to_unsigned(12443, 16)), -- 12443 / 0x309b -- last item of row
    2457 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    2458 => std_logic_vector(to_unsigned(12613, 16)), -- 12613 / 0x3145
    2459 => std_logic_vector(to_unsigned( 4431, 16)), --  4431 / 0x114f -- last item of row
    2460 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    2461 => std_logic_vector(to_unsigned( 1344, 16)), --  1344 / 0x0540
    2462 => std_logic_vector(to_unsigned( 4014, 16)), --  4014 / 0x0fae -- last item of row
    2463 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    2464 => std_logic_vector(to_unsigned( 8488, 16)), --  8488 / 0x2128
    2465 => std_logic_vector(to_unsigned(13850, 16)), -- 13850 / 0x361a -- last item of row
    2466 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    2467 => std_logic_vector(to_unsigned( 1730, 16)), --  1730 / 0x06c2
    2468 => std_logic_vector(to_unsigned(14896, 16)), -- 14896 / 0x3a30 -- last item of row
    2469 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    2470 => std_logic_vector(to_unsigned(14942, 16)), -- 14942 / 0x3a5e
    2471 => std_logic_vector(to_unsigned( 7126, 16)), --  7126 / 0x1bd6 -- last item of row
    2472 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    2473 => std_logic_vector(to_unsigned(14983, 16)), -- 14983 / 0x3a87
    2474 => std_logic_vector(to_unsigned( 8863, 16)), --  8863 / 0x229f -- last item of row
    2475 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    2476 => std_logic_vector(to_unsigned( 6578, 16)), --  6578 / 0x19b2
    2477 => std_logic_vector(to_unsigned( 8564, 16)), --  8564 / 0x2174 -- last item of row
    2478 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    2479 => std_logic_vector(to_unsigned( 4947, 16)), --  4947 / 0x1353
    2480 => std_logic_vector(to_unsigned(  396, 16)), --   396 / 0x018c -- last item of row
    2481 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    2482 => std_logic_vector(to_unsigned(  297, 16)), --   297 / 0x0129
    2483 => std_logic_vector(to_unsigned(12805, 16)), -- 12805 / 0x3205 -- last item of row
    2484 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    2485 => std_logic_vector(to_unsigned(13878, 16)), -- 13878 / 0x3636
    2486 => std_logic_vector(to_unsigned( 6692, 16)), --  6692 / 0x1a24 -- last item of row
    2487 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    2488 => std_logic_vector(to_unsigned(11857, 16)), -- 11857 / 0x2e51
    2489 => std_logic_vector(to_unsigned(11186, 16)), -- 11186 / 0x2bb2 -- last item of row
    2490 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    2491 => std_logic_vector(to_unsigned(14395, 16)), -- 14395 / 0x383b
    2492 => std_logic_vector(to_unsigned(11493, 16)), -- 11493 / 0x2ce5 -- last item of row
    2493 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    2494 => std_logic_vector(to_unsigned(16145, 16)), -- 16145 / 0x3f11
    2495 => std_logic_vector(to_unsigned(12251, 16)), -- 12251 / 0x2fdb -- last item of row
    2496 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    2497 => std_logic_vector(to_unsigned(13462, 16)), -- 13462 / 0x3496
    2498 => std_logic_vector(to_unsigned( 7428, 16)), --  7428 / 0x1d04 -- last item of row
    2499 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    2500 => std_logic_vector(to_unsigned(14526, 16)), -- 14526 / 0x38be
    2501 => std_logic_vector(to_unsigned(13119, 16)), -- 13119 / 0x333f -- last item of row
    2502 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    2503 => std_logic_vector(to_unsigned( 2535, 16)), --  2535 / 0x09e7
    2504 => std_logic_vector(to_unsigned(11243, 16)), -- 11243 / 0x2beb -- last item of row
    2505 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    2506 => std_logic_vector(to_unsigned( 6465, 16)), --  6465 / 0x1941
    2507 => std_logic_vector(to_unsigned(12690, 16)), -- 12690 / 0x3192 -- last item of row
    2508 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    2509 => std_logic_vector(to_unsigned( 6872, 16)), --  6872 / 0x1ad8
    2510 => std_logic_vector(to_unsigned( 9334, 16)), --  9334 / 0x2476 -- last item of row
    2511 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    2512 => std_logic_vector(to_unsigned(15371, 16)), -- 15371 / 0x3c0b
    2513 => std_logic_vector(to_unsigned(14023, 16)), -- 14023 / 0x36c7 -- last item of row
    2514 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    2515 => std_logic_vector(to_unsigned( 8101, 16)), --  8101 / 0x1fa5
    2516 => std_logic_vector(to_unsigned(10187, 16)), -- 10187 / 0x27cb -- last item of row
    2517 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    2518 => std_logic_vector(to_unsigned(11963, 16)), -- 11963 / 0x2ebb
    2519 => std_logic_vector(to_unsigned( 4848, 16)), --  4848 / 0x12f0 -- last item of row
    2520 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    2521 => std_logic_vector(to_unsigned(15125, 16)), -- 15125 / 0x3b15
    2522 => std_logic_vector(to_unsigned( 6119, 16)), --  6119 / 0x17e7 -- last item of row
    2523 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    2524 => std_logic_vector(to_unsigned( 8051, 16)), --  8051 / 0x1f73
    2525 => std_logic_vector(to_unsigned(14465, 16)), -- 14465 / 0x3881 -- last item of row
    2526 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    2527 => std_logic_vector(to_unsigned(11139, 16)), -- 11139 / 0x2b83
    2528 => std_logic_vector(to_unsigned( 5167, 16)), --  5167 / 0x142f -- last item of row
    2529 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    2530 => std_logic_vector(to_unsigned( 2883, 16)), --  2883 / 0x0b43
    2531 => std_logic_vector(to_unsigned(14521, 16)), -- 14521 / 0x38b9 -- last item of row
    -- Table for fecframe_normal, C3_5
    2532 => std_logic_vector(to_unsigned(22422, 16)), -- 22422 / 0x5796
    2533 => std_logic_vector(to_unsigned(10282, 16)), -- 10282 / 0x282a
    2534 => std_logic_vector(to_unsigned(11626, 16)), -- 11626 / 0x2d6a
    2535 => std_logic_vector(to_unsigned(19997, 16)), -- 19997 / 0x4e1d
    2536 => std_logic_vector(to_unsigned(11161, 16)), -- 11161 / 0x2b99
    2537 => std_logic_vector(to_unsigned( 2922, 16)), --  2922 / 0x0b6a
    2538 => std_logic_vector(to_unsigned( 3122, 16)), --  3122 / 0x0c32
    2539 => std_logic_vector(to_unsigned(   99, 16)), --    99 / 0x0063
    2540 => std_logic_vector(to_unsigned( 5625, 16)), --  5625 / 0x15f9
    2541 => std_logic_vector(to_unsigned(17064, 16)), -- 17064 / 0x42a8
    2542 => std_logic_vector(to_unsigned( 8270, 16)), --  8270 / 0x204e
    2543 => std_logic_vector(to_unsigned(  179, 16)), --   179 / 0x00b3 -- last item of row
    2544 => std_logic_vector(to_unsigned(25087, 16)), -- 25087 / 0x61ff
    2545 => std_logic_vector(to_unsigned(16218, 16)), -- 16218 / 0x3f5a
    2546 => std_logic_vector(to_unsigned(17015, 16)), -- 17015 / 0x4277
    2547 => std_logic_vector(to_unsigned(  828, 16)), --   828 / 0x033c
    2548 => std_logic_vector(to_unsigned(20041, 16)), -- 20041 / 0x4e49
    2549 => std_logic_vector(to_unsigned(25656, 16)), -- 25656 / 0x6438
    2550 => std_logic_vector(to_unsigned( 4186, 16)), --  4186 / 0x105a
    2551 => std_logic_vector(to_unsigned(11629, 16)), -- 11629 / 0x2d6d
    2552 => std_logic_vector(to_unsigned(22599, 16)), -- 22599 / 0x5847
    2553 => std_logic_vector(to_unsigned(17305, 16)), -- 17305 / 0x4399
    2554 => std_logic_vector(to_unsigned(22515, 16)), -- 22515 / 0x57f3
    2555 => std_logic_vector(to_unsigned( 6463, 16)), --  6463 / 0x193f -- last item of row
    2556 => std_logic_vector(to_unsigned(11049, 16)), -- 11049 / 0x2b29
    2557 => std_logic_vector(to_unsigned(22853, 16)), -- 22853 / 0x5945
    2558 => std_logic_vector(to_unsigned(25706, 16)), -- 25706 / 0x646a
    2559 => std_logic_vector(to_unsigned(14388, 16)), -- 14388 / 0x3834
    2560 => std_logic_vector(to_unsigned( 5500, 16)), --  5500 / 0x157c
    2561 => std_logic_vector(to_unsigned(19245, 16)), -- 19245 / 0x4b2d
    2562 => std_logic_vector(to_unsigned( 8732, 16)), --  8732 / 0x221c
    2563 => std_logic_vector(to_unsigned( 2177, 16)), --  2177 / 0x0881
    2564 => std_logic_vector(to_unsigned(13555, 16)), -- 13555 / 0x34f3
    2565 => std_logic_vector(to_unsigned(11346, 16)), -- 11346 / 0x2c52
    2566 => std_logic_vector(to_unsigned(17265, 16)), -- 17265 / 0x4371
    2567 => std_logic_vector(to_unsigned( 3069, 16)), --  3069 / 0x0bfd -- last item of row
    2568 => std_logic_vector(to_unsigned(16581, 16)), -- 16581 / 0x40c5
    2569 => std_logic_vector(to_unsigned(22225, 16)), -- 22225 / 0x56d1
    2570 => std_logic_vector(to_unsigned(12563, 16)), -- 12563 / 0x3113
    2571 => std_logic_vector(to_unsigned(19717, 16)), -- 19717 / 0x4d05
    2572 => std_logic_vector(to_unsigned(23577, 16)), -- 23577 / 0x5c19
    2573 => std_logic_vector(to_unsigned(11555, 16)), -- 11555 / 0x2d23
    2574 => std_logic_vector(to_unsigned(25496, 16)), -- 25496 / 0x6398
    2575 => std_logic_vector(to_unsigned( 6853, 16)), --  6853 / 0x1ac5
    2576 => std_logic_vector(to_unsigned(25403, 16)), -- 25403 / 0x633b
    2577 => std_logic_vector(to_unsigned( 5218, 16)), --  5218 / 0x1462
    2578 => std_logic_vector(to_unsigned(15925, 16)), -- 15925 / 0x3e35
    2579 => std_logic_vector(to_unsigned(21766, 16)), -- 21766 / 0x5506 -- last item of row
    2580 => std_logic_vector(to_unsigned(16529, 16)), -- 16529 / 0x4091
    2581 => std_logic_vector(to_unsigned(14487, 16)), -- 14487 / 0x3897
    2582 => std_logic_vector(to_unsigned( 7643, 16)), --  7643 / 0x1ddb
    2583 => std_logic_vector(to_unsigned(10715, 16)), -- 10715 / 0x29db
    2584 => std_logic_vector(to_unsigned(17442, 16)), -- 17442 / 0x4422
    2585 => std_logic_vector(to_unsigned(11119, 16)), -- 11119 / 0x2b6f
    2586 => std_logic_vector(to_unsigned( 5679, 16)), --  5679 / 0x162f
    2587 => std_logic_vector(to_unsigned(14155, 16)), -- 14155 / 0x374b
    2588 => std_logic_vector(to_unsigned(24213, 16)), -- 24213 / 0x5e95
    2589 => std_logic_vector(to_unsigned(21000, 16)), -- 21000 / 0x5208
    2590 => std_logic_vector(to_unsigned( 1116, 16)), --  1116 / 0x045c
    2591 => std_logic_vector(to_unsigned(15620, 16)), -- 15620 / 0x3d04 -- last item of row
    2592 => std_logic_vector(to_unsigned( 5340, 16)), --  5340 / 0x14dc
    2593 => std_logic_vector(to_unsigned( 8636, 16)), --  8636 / 0x21bc
    2594 => std_logic_vector(to_unsigned(16693, 16)), -- 16693 / 0x4135
    2595 => std_logic_vector(to_unsigned( 1434, 16)), --  1434 / 0x059a
    2596 => std_logic_vector(to_unsigned( 5635, 16)), --  5635 / 0x1603
    2597 => std_logic_vector(to_unsigned( 6516, 16)), --  6516 / 0x1974
    2598 => std_logic_vector(to_unsigned( 9482, 16)), --  9482 / 0x250a
    2599 => std_logic_vector(to_unsigned(20189, 16)), -- 20189 / 0x4edd
    2600 => std_logic_vector(to_unsigned( 1066, 16)), --  1066 / 0x042a
    2601 => std_logic_vector(to_unsigned(15013, 16)), -- 15013 / 0x3aa5
    2602 => std_logic_vector(to_unsigned(25361, 16)), -- 25361 / 0x6311
    2603 => std_logic_vector(to_unsigned(14243, 16)), -- 14243 / 0x37a3 -- last item of row
    2604 => std_logic_vector(to_unsigned(18506, 16)), -- 18506 / 0x484a
    2605 => std_logic_vector(to_unsigned(22236, 16)), -- 22236 / 0x56dc
    2606 => std_logic_vector(to_unsigned(20912, 16)), -- 20912 / 0x51b0
    2607 => std_logic_vector(to_unsigned( 8952, 16)), --  8952 / 0x22f8
    2608 => std_logic_vector(to_unsigned( 5421, 16)), --  5421 / 0x152d
    2609 => std_logic_vector(to_unsigned(15691, 16)), -- 15691 / 0x3d4b
    2610 => std_logic_vector(to_unsigned( 6126, 16)), --  6126 / 0x17ee
    2611 => std_logic_vector(to_unsigned(21595, 16)), -- 21595 / 0x545b
    2612 => std_logic_vector(to_unsigned(  500, 16)), --   500 / 0x01f4
    2613 => std_logic_vector(to_unsigned( 6904, 16)), --  6904 / 0x1af8
    2614 => std_logic_vector(to_unsigned(13059, 16)), -- 13059 / 0x3303
    2615 => std_logic_vector(to_unsigned( 6802, 16)), --  6802 / 0x1a92 -- last item of row
    2616 => std_logic_vector(to_unsigned( 8433, 16)), --  8433 / 0x20f1
    2617 => std_logic_vector(to_unsigned( 4694, 16)), --  4694 / 0x1256
    2618 => std_logic_vector(to_unsigned( 5524, 16)), --  5524 / 0x1594
    2619 => std_logic_vector(to_unsigned(14216, 16)), -- 14216 / 0x3788
    2620 => std_logic_vector(to_unsigned( 3685, 16)), --  3685 / 0x0e65
    2621 => std_logic_vector(to_unsigned(19721, 16)), -- 19721 / 0x4d09
    2622 => std_logic_vector(to_unsigned(25420, 16)), -- 25420 / 0x634c
    2623 => std_logic_vector(to_unsigned( 9937, 16)), --  9937 / 0x26d1
    2624 => std_logic_vector(to_unsigned(23813, 16)), -- 23813 / 0x5d05
    2625 => std_logic_vector(to_unsigned( 9047, 16)), --  9047 / 0x2357
    2626 => std_logic_vector(to_unsigned(25651, 16)), -- 25651 / 0x6433
    2627 => std_logic_vector(to_unsigned(16826, 16)), -- 16826 / 0x41ba -- last item of row
    2628 => std_logic_vector(to_unsigned(21500, 16)), -- 21500 / 0x53fc
    2629 => std_logic_vector(to_unsigned(24814, 16)), -- 24814 / 0x60ee
    2630 => std_logic_vector(to_unsigned( 6344, 16)), --  6344 / 0x18c8
    2631 => std_logic_vector(to_unsigned(17382, 16)), -- 17382 / 0x43e6
    2632 => std_logic_vector(to_unsigned( 7064, 16)), --  7064 / 0x1b98
    2633 => std_logic_vector(to_unsigned(13929, 16)), -- 13929 / 0x3669
    2634 => std_logic_vector(to_unsigned( 4004, 16)), --  4004 / 0x0fa4
    2635 => std_logic_vector(to_unsigned(16552, 16)), -- 16552 / 0x40a8
    2636 => std_logic_vector(to_unsigned(12818, 16)), -- 12818 / 0x3212
    2637 => std_logic_vector(to_unsigned( 8720, 16)), --  8720 / 0x2210
    2638 => std_logic_vector(to_unsigned( 5286, 16)), --  5286 / 0x14a6
    2639 => std_logic_vector(to_unsigned( 2206, 16)), --  2206 / 0x089e -- last item of row
    2640 => std_logic_vector(to_unsigned(22517, 16)), -- 22517 / 0x57f5
    2641 => std_logic_vector(to_unsigned( 2429, 16)), --  2429 / 0x097d
    2642 => std_logic_vector(to_unsigned(19065, 16)), -- 19065 / 0x4a79
    2643 => std_logic_vector(to_unsigned( 2921, 16)), --  2921 / 0x0b69
    2644 => std_logic_vector(to_unsigned(21611, 16)), -- 21611 / 0x546b
    2645 => std_logic_vector(to_unsigned( 1873, 16)), --  1873 / 0x0751
    2646 => std_logic_vector(to_unsigned( 7507, 16)), --  7507 / 0x1d53
    2647 => std_logic_vector(to_unsigned( 5661, 16)), --  5661 / 0x161d
    2648 => std_logic_vector(to_unsigned(23006, 16)), -- 23006 / 0x59de
    2649 => std_logic_vector(to_unsigned(23128, 16)), -- 23128 / 0x5a58
    2650 => std_logic_vector(to_unsigned(20543, 16)), -- 20543 / 0x503f
    2651 => std_logic_vector(to_unsigned(19777, 16)), -- 19777 / 0x4d41 -- last item of row
    2652 => std_logic_vector(to_unsigned( 1770, 16)), --  1770 / 0x06ea
    2653 => std_logic_vector(to_unsigned( 4636, 16)), --  4636 / 0x121c
    2654 => std_logic_vector(to_unsigned(20900, 16)), -- 20900 / 0x51a4
    2655 => std_logic_vector(to_unsigned(14931, 16)), -- 14931 / 0x3a53
    2656 => std_logic_vector(to_unsigned( 9247, 16)), --  9247 / 0x241f
    2657 => std_logic_vector(to_unsigned(12340, 16)), -- 12340 / 0x3034
    2658 => std_logic_vector(to_unsigned(11008, 16)), -- 11008 / 0x2b00
    2659 => std_logic_vector(to_unsigned(12966, 16)), -- 12966 / 0x32a6
    2660 => std_logic_vector(to_unsigned( 4471, 16)), --  4471 / 0x1177
    2661 => std_logic_vector(to_unsigned( 2731, 16)), --  2731 / 0x0aab
    2662 => std_logic_vector(to_unsigned(16445, 16)), -- 16445 / 0x403d
    2663 => std_logic_vector(to_unsigned(  791, 16)), --   791 / 0x0317 -- last item of row
    2664 => std_logic_vector(to_unsigned( 6635, 16)), --  6635 / 0x19eb
    2665 => std_logic_vector(to_unsigned(14556, 16)), -- 14556 / 0x38dc
    2666 => std_logic_vector(to_unsigned(18865, 16)), -- 18865 / 0x49b1
    2667 => std_logic_vector(to_unsigned(22421, 16)), -- 22421 / 0x5795
    2668 => std_logic_vector(to_unsigned(22124, 16)), -- 22124 / 0x566c
    2669 => std_logic_vector(to_unsigned(12697, 16)), -- 12697 / 0x3199
    2670 => std_logic_vector(to_unsigned( 9803, 16)), --  9803 / 0x264b
    2671 => std_logic_vector(to_unsigned(25485, 16)), -- 25485 / 0x638d
    2672 => std_logic_vector(to_unsigned( 7744, 16)), --  7744 / 0x1e40
    2673 => std_logic_vector(to_unsigned(18254, 16)), -- 18254 / 0x474e
    2674 => std_logic_vector(to_unsigned(11313, 16)), -- 11313 / 0x2c31
    2675 => std_logic_vector(to_unsigned( 9004, 16)), --  9004 / 0x232c -- last item of row
    2676 => std_logic_vector(to_unsigned(19982, 16)), -- 19982 / 0x4e0e
    2677 => std_logic_vector(to_unsigned(23963, 16)), -- 23963 / 0x5d9b
    2678 => std_logic_vector(to_unsigned(18912, 16)), -- 18912 / 0x49e0
    2679 => std_logic_vector(to_unsigned( 7206, 16)), --  7206 / 0x1c26
    2680 => std_logic_vector(to_unsigned(12500, 16)), -- 12500 / 0x30d4
    2681 => std_logic_vector(to_unsigned( 4382, 16)), --  4382 / 0x111e
    2682 => std_logic_vector(to_unsigned(20067, 16)), -- 20067 / 0x4e63
    2683 => std_logic_vector(to_unsigned( 6177, 16)), --  6177 / 0x1821
    2684 => std_logic_vector(to_unsigned(21007, 16)), -- 21007 / 0x520f
    2685 => std_logic_vector(to_unsigned( 1195, 16)), --  1195 / 0x04ab
    2686 => std_logic_vector(to_unsigned(23547, 16)), -- 23547 / 0x5bfb
    2687 => std_logic_vector(to_unsigned(24837, 16)), -- 24837 / 0x6105 -- last item of row
    2688 => std_logic_vector(to_unsigned(  756, 16)), --   756 / 0x02f4
    2689 => std_logic_vector(to_unsigned(11158, 16)), -- 11158 / 0x2b96
    2690 => std_logic_vector(to_unsigned(14646, 16)), -- 14646 / 0x3936
    2691 => std_logic_vector(to_unsigned(20534, 16)), -- 20534 / 0x5036
    2692 => std_logic_vector(to_unsigned( 3647, 16)), --  3647 / 0x0e3f
    2693 => std_logic_vector(to_unsigned(17728, 16)), -- 17728 / 0x4540
    2694 => std_logic_vector(to_unsigned(11676, 16)), -- 11676 / 0x2d9c
    2695 => std_logic_vector(to_unsigned(11843, 16)), -- 11843 / 0x2e43
    2696 => std_logic_vector(to_unsigned(12937, 16)), -- 12937 / 0x3289
    2697 => std_logic_vector(to_unsigned( 4402, 16)), --  4402 / 0x1132
    2698 => std_logic_vector(to_unsigned( 8261, 16)), --  8261 / 0x2045
    2699 => std_logic_vector(to_unsigned(22944, 16)), -- 22944 / 0x59a0 -- last item of row
    2700 => std_logic_vector(to_unsigned( 9306, 16)), --  9306 / 0x245a
    2701 => std_logic_vector(to_unsigned(24009, 16)), -- 24009 / 0x5dc9
    2702 => std_logic_vector(to_unsigned(10012, 16)), -- 10012 / 0x271c
    2703 => std_logic_vector(to_unsigned(11081, 16)), -- 11081 / 0x2b49
    2704 => std_logic_vector(to_unsigned( 3746, 16)), --  3746 / 0x0ea2
    2705 => std_logic_vector(to_unsigned(24325, 16)), -- 24325 / 0x5f05
    2706 => std_logic_vector(to_unsigned( 8060, 16)), --  8060 / 0x1f7c
    2707 => std_logic_vector(to_unsigned(19826, 16)), -- 19826 / 0x4d72
    2708 => std_logic_vector(to_unsigned(  842, 16)), --   842 / 0x034a
    2709 => std_logic_vector(to_unsigned( 8836, 16)), --  8836 / 0x2284
    2710 => std_logic_vector(to_unsigned( 2898, 16)), --  2898 / 0x0b52
    2711 => std_logic_vector(to_unsigned( 5019, 16)), --  5019 / 0x139b -- last item of row
    2712 => std_logic_vector(to_unsigned( 7575, 16)), --  7575 / 0x1d97
    2713 => std_logic_vector(to_unsigned( 7455, 16)), --  7455 / 0x1d1f
    2714 => std_logic_vector(to_unsigned(25244, 16)), -- 25244 / 0x629c
    2715 => std_logic_vector(to_unsigned( 4736, 16)), --  4736 / 0x1280
    2716 => std_logic_vector(to_unsigned(14400, 16)), -- 14400 / 0x3840
    2717 => std_logic_vector(to_unsigned(22981, 16)), -- 22981 / 0x59c5
    2718 => std_logic_vector(to_unsigned( 5543, 16)), --  5543 / 0x15a7
    2719 => std_logic_vector(to_unsigned( 8006, 16)), --  8006 / 0x1f46
    2720 => std_logic_vector(to_unsigned(24203, 16)), -- 24203 / 0x5e8b
    2721 => std_logic_vector(to_unsigned(13053, 16)), -- 13053 / 0x32fd
    2722 => std_logic_vector(to_unsigned( 1120, 16)), --  1120 / 0x0460
    2723 => std_logic_vector(to_unsigned( 5128, 16)), --  5128 / 0x1408 -- last item of row
    2724 => std_logic_vector(to_unsigned( 3482, 16)), --  3482 / 0x0d9a
    2725 => std_logic_vector(to_unsigned( 9270, 16)), --  9270 / 0x2436
    2726 => std_logic_vector(to_unsigned(13059, 16)), -- 13059 / 0x3303
    2727 => std_logic_vector(to_unsigned(15825, 16)), -- 15825 / 0x3dd1
    2728 => std_logic_vector(to_unsigned( 7453, 16)), --  7453 / 0x1d1d
    2729 => std_logic_vector(to_unsigned(23747, 16)), -- 23747 / 0x5cc3
    2730 => std_logic_vector(to_unsigned( 3656, 16)), --  3656 / 0x0e48
    2731 => std_logic_vector(to_unsigned(24585, 16)), -- 24585 / 0x6009
    2732 => std_logic_vector(to_unsigned(16542, 16)), -- 16542 / 0x409e
    2733 => std_logic_vector(to_unsigned(17507, 16)), -- 17507 / 0x4463
    2734 => std_logic_vector(to_unsigned(22462, 16)), -- 22462 / 0x57be
    2735 => std_logic_vector(to_unsigned(14670, 16)), -- 14670 / 0x394e -- last item of row
    2736 => std_logic_vector(to_unsigned(15627, 16)), -- 15627 / 0x3d0b
    2737 => std_logic_vector(to_unsigned(15290, 16)), -- 15290 / 0x3bba
    2738 => std_logic_vector(to_unsigned( 4198, 16)), --  4198 / 0x1066
    2739 => std_logic_vector(to_unsigned(22748, 16)), -- 22748 / 0x58dc
    2740 => std_logic_vector(to_unsigned( 5842, 16)), --  5842 / 0x16d2
    2741 => std_logic_vector(to_unsigned(13395, 16)), -- 13395 / 0x3453
    2742 => std_logic_vector(to_unsigned(23918, 16)), -- 23918 / 0x5d6e
    2743 => std_logic_vector(to_unsigned(16985, 16)), -- 16985 / 0x4259
    2744 => std_logic_vector(to_unsigned(14929, 16)), -- 14929 / 0x3a51
    2745 => std_logic_vector(to_unsigned( 3726, 16)), --  3726 / 0x0e8e
    2746 => std_logic_vector(to_unsigned(25350, 16)), -- 25350 / 0x6306
    2747 => std_logic_vector(to_unsigned(24157, 16)), -- 24157 / 0x5e5d -- last item of row
    2748 => std_logic_vector(to_unsigned(24896, 16)), -- 24896 / 0x6140
    2749 => std_logic_vector(to_unsigned(16365, 16)), -- 16365 / 0x3fed
    2750 => std_logic_vector(to_unsigned(16423, 16)), -- 16423 / 0x4027
    2751 => std_logic_vector(to_unsigned(13461, 16)), -- 13461 / 0x3495
    2752 => std_logic_vector(to_unsigned(16615, 16)), -- 16615 / 0x40e7
    2753 => std_logic_vector(to_unsigned( 8107, 16)), --  8107 / 0x1fab
    2754 => std_logic_vector(to_unsigned(24741, 16)), -- 24741 / 0x60a5
    2755 => std_logic_vector(to_unsigned( 3604, 16)), --  3604 / 0x0e14
    2756 => std_logic_vector(to_unsigned(25904, 16)), -- 25904 / 0x6530
    2757 => std_logic_vector(to_unsigned( 8716, 16)), --  8716 / 0x220c
    2758 => std_logic_vector(to_unsigned( 9604, 16)), --  9604 / 0x2584
    2759 => std_logic_vector(to_unsigned(20365, 16)), -- 20365 / 0x4f8d -- last item of row
    2760 => std_logic_vector(to_unsigned( 3729, 16)), --  3729 / 0x0e91
    2761 => std_logic_vector(to_unsigned(17245, 16)), -- 17245 / 0x435d
    2762 => std_logic_vector(to_unsigned(18448, 16)), -- 18448 / 0x4810
    2763 => std_logic_vector(to_unsigned( 9862, 16)), --  9862 / 0x2686
    2764 => std_logic_vector(to_unsigned(20831, 16)), -- 20831 / 0x515f
    2765 => std_logic_vector(to_unsigned(25326, 16)), -- 25326 / 0x62ee
    2766 => std_logic_vector(to_unsigned(20517, 16)), -- 20517 / 0x5025
    2767 => std_logic_vector(to_unsigned(24618, 16)), -- 24618 / 0x602a
    2768 => std_logic_vector(to_unsigned(13282, 16)), -- 13282 / 0x33e2
    2769 => std_logic_vector(to_unsigned( 5099, 16)), --  5099 / 0x13eb
    2770 => std_logic_vector(to_unsigned(14183, 16)), -- 14183 / 0x3767
    2771 => std_logic_vector(to_unsigned( 8804, 16)), --  8804 / 0x2264 -- last item of row
    2772 => std_logic_vector(to_unsigned(16455, 16)), -- 16455 / 0x4047
    2773 => std_logic_vector(to_unsigned(17646, 16)), -- 17646 / 0x44ee
    2774 => std_logic_vector(to_unsigned(15376, 16)), -- 15376 / 0x3c10
    2775 => std_logic_vector(to_unsigned(18194, 16)), -- 18194 / 0x4712
    2776 => std_logic_vector(to_unsigned(25528, 16)), -- 25528 / 0x63b8
    2777 => std_logic_vector(to_unsigned( 1777, 16)), --  1777 / 0x06f1
    2778 => std_logic_vector(to_unsigned( 6066, 16)), --  6066 / 0x17b2
    2779 => std_logic_vector(to_unsigned(21855, 16)), -- 21855 / 0x555f
    2780 => std_logic_vector(to_unsigned(14372, 16)), -- 14372 / 0x3824
    2781 => std_logic_vector(to_unsigned(12517, 16)), -- 12517 / 0x30e5
    2782 => std_logic_vector(to_unsigned( 4488, 16)), --  4488 / 0x1188
    2783 => std_logic_vector(to_unsigned(17490, 16)), -- 17490 / 0x4452 -- last item of row
    2784 => std_logic_vector(to_unsigned( 1400, 16)), --  1400 / 0x0578
    2785 => std_logic_vector(to_unsigned( 8135, 16)), --  8135 / 0x1fc7
    2786 => std_logic_vector(to_unsigned(23375, 16)), -- 23375 / 0x5b4f
    2787 => std_logic_vector(to_unsigned(20879, 16)), -- 20879 / 0x518f
    2788 => std_logic_vector(to_unsigned( 8476, 16)), --  8476 / 0x211c
    2789 => std_logic_vector(to_unsigned( 4084, 16)), --  4084 / 0x0ff4
    2790 => std_logic_vector(to_unsigned(12936, 16)), -- 12936 / 0x3288
    2791 => std_logic_vector(to_unsigned(25536, 16)), -- 25536 / 0x63c0
    2792 => std_logic_vector(to_unsigned(22309, 16)), -- 22309 / 0x5725
    2793 => std_logic_vector(to_unsigned(16582, 16)), -- 16582 / 0x40c6
    2794 => std_logic_vector(to_unsigned( 6402, 16)), --  6402 / 0x1902
    2795 => std_logic_vector(to_unsigned(24360, 16)), -- 24360 / 0x5f28 -- last item of row
    2796 => std_logic_vector(to_unsigned(25119, 16)), -- 25119 / 0x621f
    2797 => std_logic_vector(to_unsigned(23586, 16)), -- 23586 / 0x5c22
    2798 => std_logic_vector(to_unsigned(  128, 16)), --   128 / 0x0080
    2799 => std_logic_vector(to_unsigned( 4761, 16)), --  4761 / 0x1299
    2800 => std_logic_vector(to_unsigned(10443, 16)), -- 10443 / 0x28cb
    2801 => std_logic_vector(to_unsigned(22536, 16)), -- 22536 / 0x5808
    2802 => std_logic_vector(to_unsigned( 8607, 16)), --  8607 / 0x219f
    2803 => std_logic_vector(to_unsigned( 9752, 16)), --  9752 / 0x2618
    2804 => std_logic_vector(to_unsigned(25446, 16)), -- 25446 / 0x6366
    2805 => std_logic_vector(to_unsigned(15053, 16)), -- 15053 / 0x3acd
    2806 => std_logic_vector(to_unsigned( 1856, 16)), --  1856 / 0x0740
    2807 => std_logic_vector(to_unsigned( 4040, 16)), --  4040 / 0x0fc8 -- last item of row
    2808 => std_logic_vector(to_unsigned(  377, 16)), --   377 / 0x0179
    2809 => std_logic_vector(to_unsigned(21160, 16)), -- 21160 / 0x52a8
    2810 => std_logic_vector(to_unsigned(13474, 16)), -- 13474 / 0x34a2
    2811 => std_logic_vector(to_unsigned( 5451, 16)), --  5451 / 0x154b
    2812 => std_logic_vector(to_unsigned(17170, 16)), -- 17170 / 0x4312
    2813 => std_logic_vector(to_unsigned( 5938, 16)), --  5938 / 0x1732
    2814 => std_logic_vector(to_unsigned(10256, 16)), -- 10256 / 0x2810
    2815 => std_logic_vector(to_unsigned(11972, 16)), -- 11972 / 0x2ec4
    2816 => std_logic_vector(to_unsigned(24210, 16)), -- 24210 / 0x5e92
    2817 => std_logic_vector(to_unsigned(17833, 16)), -- 17833 / 0x45a9
    2818 => std_logic_vector(to_unsigned(22047, 16)), -- 22047 / 0x561f
    2819 => std_logic_vector(to_unsigned(16108, 16)), -- 16108 / 0x3eec -- last item of row
    2820 => std_logic_vector(to_unsigned(13075, 16)), -- 13075 / 0x3313
    2821 => std_logic_vector(to_unsigned( 9648, 16)), --  9648 / 0x25b0
    2822 => std_logic_vector(to_unsigned(24546, 16)), -- 24546 / 0x5fe2
    2823 => std_logic_vector(to_unsigned(13150, 16)), -- 13150 / 0x335e
    2824 => std_logic_vector(to_unsigned(23867, 16)), -- 23867 / 0x5d3b
    2825 => std_logic_vector(to_unsigned( 7309, 16)), --  7309 / 0x1c8d
    2826 => std_logic_vector(to_unsigned(19798, 16)), -- 19798 / 0x4d56
    2827 => std_logic_vector(to_unsigned( 2988, 16)), --  2988 / 0x0bac
    2828 => std_logic_vector(to_unsigned(16858, 16)), -- 16858 / 0x41da
    2829 => std_logic_vector(to_unsigned( 4825, 16)), --  4825 / 0x12d9
    2830 => std_logic_vector(to_unsigned(23950, 16)), -- 23950 / 0x5d8e
    2831 => std_logic_vector(to_unsigned(15125, 16)), -- 15125 / 0x3b15 -- last item of row
    2832 => std_logic_vector(to_unsigned(20526, 16)), -- 20526 / 0x502e
    2833 => std_logic_vector(to_unsigned( 3553, 16)), --  3553 / 0x0de1
    2834 => std_logic_vector(to_unsigned(11525, 16)), -- 11525 / 0x2d05
    2835 => std_logic_vector(to_unsigned(23366, 16)), -- 23366 / 0x5b46
    2836 => std_logic_vector(to_unsigned( 2452, 16)), --  2452 / 0x0994
    2837 => std_logic_vector(to_unsigned(17626, 16)), -- 17626 / 0x44da
    2838 => std_logic_vector(to_unsigned(19265, 16)), -- 19265 / 0x4b41
    2839 => std_logic_vector(to_unsigned(20172, 16)), -- 20172 / 0x4ecc
    2840 => std_logic_vector(to_unsigned(18060, 16)), -- 18060 / 0x468c
    2841 => std_logic_vector(to_unsigned(24593, 16)), -- 24593 / 0x6011
    2842 => std_logic_vector(to_unsigned(13255, 16)), -- 13255 / 0x33c7
    2843 => std_logic_vector(to_unsigned( 1552, 16)), --  1552 / 0x0610 -- last item of row
    2844 => std_logic_vector(to_unsigned(18839, 16)), -- 18839 / 0x4997
    2845 => std_logic_vector(to_unsigned(21132, 16)), -- 21132 / 0x528c
    2846 => std_logic_vector(to_unsigned(20119, 16)), -- 20119 / 0x4e97
    2847 => std_logic_vector(to_unsigned(15214, 16)), -- 15214 / 0x3b6e
    2848 => std_logic_vector(to_unsigned(14705, 16)), -- 14705 / 0x3971
    2849 => std_logic_vector(to_unsigned( 7096, 16)), --  7096 / 0x1bb8
    2850 => std_logic_vector(to_unsigned(10174, 16)), -- 10174 / 0x27be
    2851 => std_logic_vector(to_unsigned( 5663, 16)), --  5663 / 0x161f
    2852 => std_logic_vector(to_unsigned(18651, 16)), -- 18651 / 0x48db
    2853 => std_logic_vector(to_unsigned(19700, 16)), -- 19700 / 0x4cf4
    2854 => std_logic_vector(to_unsigned(12524, 16)), -- 12524 / 0x30ec
    2855 => std_logic_vector(to_unsigned(14033, 16)), -- 14033 / 0x36d1 -- last item of row
    2856 => std_logic_vector(to_unsigned( 4127, 16)), --  4127 / 0x101f
    2857 => std_logic_vector(to_unsigned( 2971, 16)), --  2971 / 0x0b9b
    2858 => std_logic_vector(to_unsigned(17499, 16)), -- 17499 / 0x445b
    2859 => std_logic_vector(to_unsigned(16287, 16)), -- 16287 / 0x3f9f
    2860 => std_logic_vector(to_unsigned(22368, 16)), -- 22368 / 0x5760
    2861 => std_logic_vector(to_unsigned(21463, 16)), -- 21463 / 0x53d7
    2862 => std_logic_vector(to_unsigned( 7943, 16)), --  7943 / 0x1f07
    2863 => std_logic_vector(to_unsigned(18880, 16)), -- 18880 / 0x49c0
    2864 => std_logic_vector(to_unsigned( 5567, 16)), --  5567 / 0x15bf
    2865 => std_logic_vector(to_unsigned( 8047, 16)), --  8047 / 0x1f6f
    2866 => std_logic_vector(to_unsigned(23363, 16)), -- 23363 / 0x5b43
    2867 => std_logic_vector(to_unsigned( 6797, 16)), --  6797 / 0x1a8d -- last item of row
    2868 => std_logic_vector(to_unsigned(10651, 16)), -- 10651 / 0x299b
    2869 => std_logic_vector(to_unsigned(24471, 16)), -- 24471 / 0x5f97
    2870 => std_logic_vector(to_unsigned(14325, 16)), -- 14325 / 0x37f5
    2871 => std_logic_vector(to_unsigned( 4081, 16)), --  4081 / 0x0ff1
    2872 => std_logic_vector(to_unsigned( 7258, 16)), --  7258 / 0x1c5a
    2873 => std_logic_vector(to_unsigned( 4949, 16)), --  4949 / 0x1355
    2874 => std_logic_vector(to_unsigned( 7044, 16)), --  7044 / 0x1b84
    2875 => std_logic_vector(to_unsigned( 1078, 16)), --  1078 / 0x0436
    2876 => std_logic_vector(to_unsigned(  797, 16)), --   797 / 0x031d
    2877 => std_logic_vector(to_unsigned(22910, 16)), -- 22910 / 0x597e
    2878 => std_logic_vector(to_unsigned(20474, 16)), -- 20474 / 0x4ffa
    2879 => std_logic_vector(to_unsigned( 4318, 16)), --  4318 / 0x10de -- last item of row
    2880 => std_logic_vector(to_unsigned(21374, 16)), -- 21374 / 0x537e
    2881 => std_logic_vector(to_unsigned(13231, 16)), -- 13231 / 0x33af
    2882 => std_logic_vector(to_unsigned(22985, 16)), -- 22985 / 0x59c9
    2883 => std_logic_vector(to_unsigned( 5056, 16)), --  5056 / 0x13c0
    2884 => std_logic_vector(to_unsigned( 3821, 16)), --  3821 / 0x0eed
    2885 => std_logic_vector(to_unsigned(23718, 16)), -- 23718 / 0x5ca6
    2886 => std_logic_vector(to_unsigned(14178, 16)), -- 14178 / 0x3762
    2887 => std_logic_vector(to_unsigned( 9978, 16)), --  9978 / 0x26fa
    2888 => std_logic_vector(to_unsigned(19030, 16)), -- 19030 / 0x4a56
    2889 => std_logic_vector(to_unsigned(23594, 16)), -- 23594 / 0x5c2a
    2890 => std_logic_vector(to_unsigned( 8895, 16)), --  8895 / 0x22bf
    2891 => std_logic_vector(to_unsigned(25358, 16)), -- 25358 / 0x630e -- last item of row
    2892 => std_logic_vector(to_unsigned( 6199, 16)), --  6199 / 0x1837
    2893 => std_logic_vector(to_unsigned(22056, 16)), -- 22056 / 0x5628
    2894 => std_logic_vector(to_unsigned( 7749, 16)), --  7749 / 0x1e45
    2895 => std_logic_vector(to_unsigned(13310, 16)), -- 13310 / 0x33fe
    2896 => std_logic_vector(to_unsigned( 3999, 16)), --  3999 / 0x0f9f
    2897 => std_logic_vector(to_unsigned(23697, 16)), -- 23697 / 0x5c91
    2898 => std_logic_vector(to_unsigned(16445, 16)), -- 16445 / 0x403d
    2899 => std_logic_vector(to_unsigned(22636, 16)), -- 22636 / 0x586c
    2900 => std_logic_vector(to_unsigned( 5225, 16)), --  5225 / 0x1469
    2901 => std_logic_vector(to_unsigned(22437, 16)), -- 22437 / 0x57a5
    2902 => std_logic_vector(to_unsigned(24153, 16)), -- 24153 / 0x5e59
    2903 => std_logic_vector(to_unsigned( 9442, 16)), --  9442 / 0x24e2 -- last item of row
    2904 => std_logic_vector(to_unsigned( 7978, 16)), --  7978 / 0x1f2a
    2905 => std_logic_vector(to_unsigned(12177, 16)), -- 12177 / 0x2f91
    2906 => std_logic_vector(to_unsigned( 2893, 16)), --  2893 / 0x0b4d
    2907 => std_logic_vector(to_unsigned(20778, 16)), -- 20778 / 0x512a
    2908 => std_logic_vector(to_unsigned( 3175, 16)), --  3175 / 0x0c67
    2909 => std_logic_vector(to_unsigned( 8645, 16)), --  8645 / 0x21c5
    2910 => std_logic_vector(to_unsigned(11863, 16)), -- 11863 / 0x2e57
    2911 => std_logic_vector(to_unsigned(24623, 16)), -- 24623 / 0x602f
    2912 => std_logic_vector(to_unsigned(10311, 16)), -- 10311 / 0x2847
    2913 => std_logic_vector(to_unsigned(25767, 16)), -- 25767 / 0x64a7
    2914 => std_logic_vector(to_unsigned(17057, 16)), -- 17057 / 0x42a1
    2915 => std_logic_vector(to_unsigned( 3691, 16)), --  3691 / 0x0e6b -- last item of row
    2916 => std_logic_vector(to_unsigned(20473, 16)), -- 20473 / 0x4ff9
    2917 => std_logic_vector(to_unsigned(11294, 16)), -- 11294 / 0x2c1e
    2918 => std_logic_vector(to_unsigned( 9914, 16)), --  9914 / 0x26ba
    2919 => std_logic_vector(to_unsigned(22815, 16)), -- 22815 / 0x591f
    2920 => std_logic_vector(to_unsigned( 2574, 16)), --  2574 / 0x0a0e
    2921 => std_logic_vector(to_unsigned( 8439, 16)), --  8439 / 0x20f7
    2922 => std_logic_vector(to_unsigned( 3699, 16)), --  3699 / 0x0e73
    2923 => std_logic_vector(to_unsigned( 5431, 16)), --  5431 / 0x1537
    2924 => std_logic_vector(to_unsigned(24840, 16)), -- 24840 / 0x6108
    2925 => std_logic_vector(to_unsigned(21908, 16)), -- 21908 / 0x5594
    2926 => std_logic_vector(to_unsigned(16088, 16)), -- 16088 / 0x3ed8
    2927 => std_logic_vector(to_unsigned(18244, 16)), -- 18244 / 0x4744 -- last item of row
    2928 => std_logic_vector(to_unsigned( 8208, 16)), --  8208 / 0x2010
    2929 => std_logic_vector(to_unsigned( 5755, 16)), --  5755 / 0x167b
    2930 => std_logic_vector(to_unsigned(19059, 16)), -- 19059 / 0x4a73
    2931 => std_logic_vector(to_unsigned( 8541, 16)), --  8541 / 0x215d
    2932 => std_logic_vector(to_unsigned(24924, 16)), -- 24924 / 0x615c
    2933 => std_logic_vector(to_unsigned( 6454, 16)), --  6454 / 0x1936
    2934 => std_logic_vector(to_unsigned(11234, 16)), -- 11234 / 0x2be2
    2935 => std_logic_vector(to_unsigned(10492, 16)), -- 10492 / 0x28fc
    2936 => std_logic_vector(to_unsigned(16406, 16)), -- 16406 / 0x4016
    2937 => std_logic_vector(to_unsigned(10831, 16)), -- 10831 / 0x2a4f
    2938 => std_logic_vector(to_unsigned(11436, 16)), -- 11436 / 0x2cac
    2939 => std_logic_vector(to_unsigned( 9649, 16)), --  9649 / 0x25b1 -- last item of row
    2940 => std_logic_vector(to_unsigned(16264, 16)), -- 16264 / 0x3f88
    2941 => std_logic_vector(to_unsigned(11275, 16)), -- 11275 / 0x2c0b
    2942 => std_logic_vector(to_unsigned(24953, 16)), -- 24953 / 0x6179
    2943 => std_logic_vector(to_unsigned( 2347, 16)), --  2347 / 0x092b
    2944 => std_logic_vector(to_unsigned(12667, 16)), -- 12667 / 0x317b
    2945 => std_logic_vector(to_unsigned(19190, 16)), -- 19190 / 0x4af6
    2946 => std_logic_vector(to_unsigned( 7257, 16)), --  7257 / 0x1c59
    2947 => std_logic_vector(to_unsigned( 7174, 16)), --  7174 / 0x1c06
    2948 => std_logic_vector(to_unsigned(24819, 16)), -- 24819 / 0x60f3
    2949 => std_logic_vector(to_unsigned( 2938, 16)), --  2938 / 0x0b7a
    2950 => std_logic_vector(to_unsigned( 2522, 16)), --  2522 / 0x09da
    2951 => std_logic_vector(to_unsigned(11749, 16)), -- 11749 / 0x2de5 -- last item of row
    2952 => std_logic_vector(to_unsigned( 3627, 16)), --  3627 / 0x0e2b
    2953 => std_logic_vector(to_unsigned( 5969, 16)), --  5969 / 0x1751
    2954 => std_logic_vector(to_unsigned(13862, 16)), -- 13862 / 0x3626
    2955 => std_logic_vector(to_unsigned( 1538, 16)), --  1538 / 0x0602
    2956 => std_logic_vector(to_unsigned(23176, 16)), -- 23176 / 0x5a88
    2957 => std_logic_vector(to_unsigned( 6353, 16)), --  6353 / 0x18d1
    2958 => std_logic_vector(to_unsigned( 2855, 16)), --  2855 / 0x0b27
    2959 => std_logic_vector(to_unsigned(17720, 16)), -- 17720 / 0x4538
    2960 => std_logic_vector(to_unsigned( 2472, 16)), --  2472 / 0x09a8
    2961 => std_logic_vector(to_unsigned( 7428, 16)), --  7428 / 0x1d04
    2962 => std_logic_vector(to_unsigned(  573, 16)), --   573 / 0x023d
    2963 => std_logic_vector(to_unsigned(15036, 16)), -- 15036 / 0x3abc -- last item of row
    2964 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    2965 => std_logic_vector(to_unsigned(18539, 16)), -- 18539 / 0x486b
    2966 => std_logic_vector(to_unsigned(18661, 16)), -- 18661 / 0x48e5 -- last item of row
    2967 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    2968 => std_logic_vector(to_unsigned(10502, 16)), -- 10502 / 0x2906
    2969 => std_logic_vector(to_unsigned( 3002, 16)), --  3002 / 0x0bba -- last item of row
    2970 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    2971 => std_logic_vector(to_unsigned( 9368, 16)), --  9368 / 0x2498
    2972 => std_logic_vector(to_unsigned(10761, 16)), -- 10761 / 0x2a09 -- last item of row
    2973 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    2974 => std_logic_vector(to_unsigned(12299, 16)), -- 12299 / 0x300b
    2975 => std_logic_vector(to_unsigned( 7828, 16)), --  7828 / 0x1e94 -- last item of row
    2976 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    2977 => std_logic_vector(to_unsigned(15048, 16)), -- 15048 / 0x3ac8
    2978 => std_logic_vector(to_unsigned(13362, 16)), -- 13362 / 0x3432 -- last item of row
    2979 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    2980 => std_logic_vector(to_unsigned(18444, 16)), -- 18444 / 0x480c
    2981 => std_logic_vector(to_unsigned(24640, 16)), -- 24640 / 0x6040 -- last item of row
    2982 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    2983 => std_logic_vector(to_unsigned(20775, 16)), -- 20775 / 0x5127
    2984 => std_logic_vector(to_unsigned(19175, 16)), -- 19175 / 0x4ae7 -- last item of row
    2985 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    2986 => std_logic_vector(to_unsigned(18970, 16)), -- 18970 / 0x4a1a
    2987 => std_logic_vector(to_unsigned(10971, 16)), -- 10971 / 0x2adb -- last item of row
    2988 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    2989 => std_logic_vector(to_unsigned( 5329, 16)), --  5329 / 0x14d1
    2990 => std_logic_vector(to_unsigned(19982, 16)), -- 19982 / 0x4e0e -- last item of row
    2991 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    2992 => std_logic_vector(to_unsigned(11296, 16)), -- 11296 / 0x2c20
    2993 => std_logic_vector(to_unsigned(18655, 16)), -- 18655 / 0x48df -- last item of row
    2994 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    2995 => std_logic_vector(to_unsigned(15046, 16)), -- 15046 / 0x3ac6
    2996 => std_logic_vector(to_unsigned(20659, 16)), -- 20659 / 0x50b3 -- last item of row
    2997 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    2998 => std_logic_vector(to_unsigned( 7300, 16)), --  7300 / 0x1c84
    2999 => std_logic_vector(to_unsigned(22140, 16)), -- 22140 / 0x567c -- last item of row
    3000 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3001 => std_logic_vector(to_unsigned(22029, 16)), -- 22029 / 0x560d
    3002 => std_logic_vector(to_unsigned(14477, 16)), -- 14477 / 0x388d -- last item of row
    3003 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3004 => std_logic_vector(to_unsigned(11129, 16)), -- 11129 / 0x2b79
    3005 => std_logic_vector(to_unsigned(  742, 16)), --   742 / 0x02e6 -- last item of row
    3006 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3007 => std_logic_vector(to_unsigned(13254, 16)), -- 13254 / 0x33c6
    3008 => std_logic_vector(to_unsigned(13813, 16)), -- 13813 / 0x35f5 -- last item of row
    3009 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3010 => std_logic_vector(to_unsigned(19234, 16)), -- 19234 / 0x4b22
    3011 => std_logic_vector(to_unsigned(13273, 16)), -- 13273 / 0x33d9 -- last item of row
    3012 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3013 => std_logic_vector(to_unsigned( 6079, 16)), --  6079 / 0x17bf
    3014 => std_logic_vector(to_unsigned(21122, 16)), -- 21122 / 0x5282 -- last item of row
    3015 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3016 => std_logic_vector(to_unsigned(22782, 16)), -- 22782 / 0x58fe
    3017 => std_logic_vector(to_unsigned( 5828, 16)), --  5828 / 0x16c4 -- last item of row
    3018 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3019 => std_logic_vector(to_unsigned(19775, 16)), -- 19775 / 0x4d3f
    3020 => std_logic_vector(to_unsigned( 4247, 16)), --  4247 / 0x1097 -- last item of row
    3021 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3022 => std_logic_vector(to_unsigned( 1660, 16)), --  1660 / 0x067c
    3023 => std_logic_vector(to_unsigned(19413, 16)), -- 19413 / 0x4bd5 -- last item of row
    3024 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3025 => std_logic_vector(to_unsigned( 4403, 16)), --  4403 / 0x1133
    3026 => std_logic_vector(to_unsigned( 3649, 16)), --  3649 / 0x0e41 -- last item of row
    3027 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3028 => std_logic_vector(to_unsigned(13371, 16)), -- 13371 / 0x343b
    3029 => std_logic_vector(to_unsigned(25851, 16)), -- 25851 / 0x64fb -- last item of row
    3030 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3031 => std_logic_vector(to_unsigned(22770, 16)), -- 22770 / 0x58f2
    3032 => std_logic_vector(to_unsigned(21784, 16)), -- 21784 / 0x5518 -- last item of row
    3033 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3034 => std_logic_vector(to_unsigned(10757, 16)), -- 10757 / 0x2a05
    3035 => std_logic_vector(to_unsigned(14131, 16)), -- 14131 / 0x3733 -- last item of row
    3036 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3037 => std_logic_vector(to_unsigned(16071, 16)), -- 16071 / 0x3ec7
    3038 => std_logic_vector(to_unsigned(21617, 16)), -- 21617 / 0x5471 -- last item of row
    3039 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3040 => std_logic_vector(to_unsigned( 6393, 16)), --  6393 / 0x18f9
    3041 => std_logic_vector(to_unsigned( 3725, 16)), --  3725 / 0x0e8d -- last item of row
    3042 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3043 => std_logic_vector(to_unsigned(  597, 16)), --   597 / 0x0255
    3044 => std_logic_vector(to_unsigned(19968, 16)), -- 19968 / 0x4e00 -- last item of row
    3045 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3046 => std_logic_vector(to_unsigned( 5743, 16)), --  5743 / 0x166f
    3047 => std_logic_vector(to_unsigned( 8084, 16)), --  8084 / 0x1f94 -- last item of row
    3048 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3049 => std_logic_vector(to_unsigned( 6770, 16)), --  6770 / 0x1a72
    3050 => std_logic_vector(to_unsigned( 9548, 16)), --  9548 / 0x254c -- last item of row
    3051 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3052 => std_logic_vector(to_unsigned( 4285, 16)), --  4285 / 0x10bd
    3053 => std_logic_vector(to_unsigned(17542, 16)), -- 17542 / 0x4486 -- last item of row
    3054 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    3055 => std_logic_vector(to_unsigned(13568, 16)), -- 13568 / 0x3500
    3056 => std_logic_vector(to_unsigned(22599, 16)), -- 22599 / 0x5847 -- last item of row
    3057 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    3058 => std_logic_vector(to_unsigned( 1786, 16)), --  1786 / 0x06fa
    3059 => std_logic_vector(to_unsigned( 4617, 16)), --  4617 / 0x1209 -- last item of row
    3060 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    3061 => std_logic_vector(to_unsigned(23238, 16)), -- 23238 / 0x5ac6
    3062 => std_logic_vector(to_unsigned(11648, 16)), -- 11648 / 0x2d80 -- last item of row
    3063 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    3064 => std_logic_vector(to_unsigned(19627, 16)), -- 19627 / 0x4cab
    3065 => std_logic_vector(to_unsigned( 2030, 16)), --  2030 / 0x07ee -- last item of row
    3066 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    3067 => std_logic_vector(to_unsigned(13601, 16)), -- 13601 / 0x3521
    3068 => std_logic_vector(to_unsigned(13458, 16)), -- 13458 / 0x3492 -- last item of row
    3069 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    3070 => std_logic_vector(to_unsigned(13740, 16)), -- 13740 / 0x35ac
    3071 => std_logic_vector(to_unsigned(17328, 16)), -- 17328 / 0x43b0 -- last item of row
    3072 => std_logic_vector(to_unsigned(   36, 16)), --    36 / 0x0024
    3073 => std_logic_vector(to_unsigned(25012, 16)), -- 25012 / 0x61b4
    3074 => std_logic_vector(to_unsigned(13944, 16)), -- 13944 / 0x3678 -- last item of row
    3075 => std_logic_vector(to_unsigned(   37, 16)), --    37 / 0x0025
    3076 => std_logic_vector(to_unsigned(22513, 16)), -- 22513 / 0x57f1
    3077 => std_logic_vector(to_unsigned( 6687, 16)), --  6687 / 0x1a1f -- last item of row
    3078 => std_logic_vector(to_unsigned(   38, 16)), --    38 / 0x0026
    3079 => std_logic_vector(to_unsigned( 4934, 16)), --  4934 / 0x1346
    3080 => std_logic_vector(to_unsigned(12587, 16)), -- 12587 / 0x312b -- last item of row
    3081 => std_logic_vector(to_unsigned(   39, 16)), --    39 / 0x0027
    3082 => std_logic_vector(to_unsigned(21197, 16)), -- 21197 / 0x52cd
    3083 => std_logic_vector(to_unsigned( 5133, 16)), --  5133 / 0x140d -- last item of row
    3084 => std_logic_vector(to_unsigned(   40, 16)), --    40 / 0x0028
    3085 => std_logic_vector(to_unsigned(22705, 16)), -- 22705 / 0x58b1
    3086 => std_logic_vector(to_unsigned( 6938, 16)), --  6938 / 0x1b1a -- last item of row
    3087 => std_logic_vector(to_unsigned(   41, 16)), --    41 / 0x0029
    3088 => std_logic_vector(to_unsigned( 7534, 16)), --  7534 / 0x1d6e
    3089 => std_logic_vector(to_unsigned(24633, 16)), -- 24633 / 0x6039 -- last item of row
    3090 => std_logic_vector(to_unsigned(   42, 16)), --    42 / 0x002a
    3091 => std_logic_vector(to_unsigned(24400, 16)), -- 24400 / 0x5f50
    3092 => std_logic_vector(to_unsigned(12797, 16)), -- 12797 / 0x31fd -- last item of row
    3093 => std_logic_vector(to_unsigned(   43, 16)), --    43 / 0x002b
    3094 => std_logic_vector(to_unsigned(21911, 16)), -- 21911 / 0x5597
    3095 => std_logic_vector(to_unsigned(25712, 16)), -- 25712 / 0x6470 -- last item of row
    3096 => std_logic_vector(to_unsigned(   44, 16)), --    44 / 0x002c
    3097 => std_logic_vector(to_unsigned(12039, 16)), -- 12039 / 0x2f07
    3098 => std_logic_vector(to_unsigned( 1140, 16)), --  1140 / 0x0474 -- last item of row
    3099 => std_logic_vector(to_unsigned(   45, 16)), --    45 / 0x002d
    3100 => std_logic_vector(to_unsigned(24306, 16)), -- 24306 / 0x5ef2
    3101 => std_logic_vector(to_unsigned( 1021, 16)), --  1021 / 0x03fd -- last item of row
    3102 => std_logic_vector(to_unsigned(   46, 16)), --    46 / 0x002e
    3103 => std_logic_vector(to_unsigned(14012, 16)), -- 14012 / 0x36bc
    3104 => std_logic_vector(to_unsigned(20747, 16)), -- 20747 / 0x510b -- last item of row
    3105 => std_logic_vector(to_unsigned(   47, 16)), --    47 / 0x002f
    3106 => std_logic_vector(to_unsigned(11265, 16)), -- 11265 / 0x2c01
    3107 => std_logic_vector(to_unsigned(15219, 16)), -- 15219 / 0x3b73 -- last item of row
    3108 => std_logic_vector(to_unsigned(   48, 16)), --    48 / 0x0030
    3109 => std_logic_vector(to_unsigned( 4670, 16)), --  4670 / 0x123e
    3110 => std_logic_vector(to_unsigned(15531, 16)), -- 15531 / 0x3cab -- last item of row
    3111 => std_logic_vector(to_unsigned(   49, 16)), --    49 / 0x0031
    3112 => std_logic_vector(to_unsigned( 9417, 16)), --  9417 / 0x24c9
    3113 => std_logic_vector(to_unsigned(14359, 16)), -- 14359 / 0x3817 -- last item of row
    3114 => std_logic_vector(to_unsigned(   50, 16)), --    50 / 0x0032
    3115 => std_logic_vector(to_unsigned( 2415, 16)), --  2415 / 0x096f
    3116 => std_logic_vector(to_unsigned( 6504, 16)), --  6504 / 0x1968 -- last item of row
    3117 => std_logic_vector(to_unsigned(   51, 16)), --    51 / 0x0033
    3118 => std_logic_vector(to_unsigned(24964, 16)), -- 24964 / 0x6184
    3119 => std_logic_vector(to_unsigned(24690, 16)), -- 24690 / 0x6072 -- last item of row
    3120 => std_logic_vector(to_unsigned(   52, 16)), --    52 / 0x0034
    3121 => std_logic_vector(to_unsigned(14443, 16)), -- 14443 / 0x386b
    3122 => std_logic_vector(to_unsigned( 8816, 16)), --  8816 / 0x2270 -- last item of row
    3123 => std_logic_vector(to_unsigned(   53, 16)), --    53 / 0x0035
    3124 => std_logic_vector(to_unsigned( 6926, 16)), --  6926 / 0x1b0e
    3125 => std_logic_vector(to_unsigned( 1291, 16)), --  1291 / 0x050b -- last item of row
    3126 => std_logic_vector(to_unsigned(   54, 16)), --    54 / 0x0036
    3127 => std_logic_vector(to_unsigned( 6209, 16)), --  6209 / 0x1841
    3128 => std_logic_vector(to_unsigned(20806, 16)), -- 20806 / 0x5146 -- last item of row
    3129 => std_logic_vector(to_unsigned(   55, 16)), --    55 / 0x0037
    3130 => std_logic_vector(to_unsigned(13915, 16)), -- 13915 / 0x365b
    3131 => std_logic_vector(to_unsigned( 4079, 16)), --  4079 / 0x0fef -- last item of row
    3132 => std_logic_vector(to_unsigned(   56, 16)), --    56 / 0x0038
    3133 => std_logic_vector(to_unsigned(24410, 16)), -- 24410 / 0x5f5a
    3134 => std_logic_vector(to_unsigned(13196, 16)), -- 13196 / 0x338c -- last item of row
    3135 => std_logic_vector(to_unsigned(   57, 16)), --    57 / 0x0039
    3136 => std_logic_vector(to_unsigned(13505, 16)), -- 13505 / 0x34c1
    3137 => std_logic_vector(to_unsigned( 6117, 16)), --  6117 / 0x17e5 -- last item of row
    3138 => std_logic_vector(to_unsigned(   58, 16)), --    58 / 0x003a
    3139 => std_logic_vector(to_unsigned( 9869, 16)), --  9869 / 0x268d
    3140 => std_logic_vector(to_unsigned( 8220, 16)), --  8220 / 0x201c -- last item of row
    3141 => std_logic_vector(to_unsigned(   59, 16)), --    59 / 0x003b
    3142 => std_logic_vector(to_unsigned( 1570, 16)), --  1570 / 0x0622
    3143 => std_logic_vector(to_unsigned( 6044, 16)), --  6044 / 0x179c -- last item of row
    3144 => std_logic_vector(to_unsigned(   60, 16)), --    60 / 0x003c
    3145 => std_logic_vector(to_unsigned(25780, 16)), -- 25780 / 0x64b4
    3146 => std_logic_vector(to_unsigned(17387, 16)), -- 17387 / 0x43eb -- last item of row
    3147 => std_logic_vector(to_unsigned(   61, 16)), --    61 / 0x003d
    3148 => std_logic_vector(to_unsigned(20671, 16)), -- 20671 / 0x50bf
    3149 => std_logic_vector(to_unsigned(24913, 16)), -- 24913 / 0x6151 -- last item of row
    3150 => std_logic_vector(to_unsigned(   62, 16)), --    62 / 0x003e
    3151 => std_logic_vector(to_unsigned(24558, 16)), -- 24558 / 0x5fee
    3152 => std_logic_vector(to_unsigned(20591, 16)), -- 20591 / 0x506f -- last item of row
    3153 => std_logic_vector(to_unsigned(   63, 16)), --    63 / 0x003f
    3154 => std_logic_vector(to_unsigned(12402, 16)), -- 12402 / 0x3072
    3155 => std_logic_vector(to_unsigned( 3702, 16)), --  3702 / 0x0e76 -- last item of row
    3156 => std_logic_vector(to_unsigned(   64, 16)), --    64 / 0x0040
    3157 => std_logic_vector(to_unsigned( 8314, 16)), --  8314 / 0x207a
    3158 => std_logic_vector(to_unsigned( 1357, 16)), --  1357 / 0x054d -- last item of row
    3159 => std_logic_vector(to_unsigned(   65, 16)), --    65 / 0x0041
    3160 => std_logic_vector(to_unsigned(20071, 16)), -- 20071 / 0x4e67
    3161 => std_logic_vector(to_unsigned(14616, 16)), -- 14616 / 0x3918 -- last item of row
    3162 => std_logic_vector(to_unsigned(   66, 16)), --    66 / 0x0042
    3163 => std_logic_vector(to_unsigned(17014, 16)), -- 17014 / 0x4276
    3164 => std_logic_vector(to_unsigned( 3688, 16)), --  3688 / 0x0e68 -- last item of row
    3165 => std_logic_vector(to_unsigned(   67, 16)), --    67 / 0x0043
    3166 => std_logic_vector(to_unsigned(19837, 16)), -- 19837 / 0x4d7d
    3167 => std_logic_vector(to_unsigned(  946, 16)), --   946 / 0x03b2 -- last item of row
    3168 => std_logic_vector(to_unsigned(   68, 16)), --    68 / 0x0044
    3169 => std_logic_vector(to_unsigned(15195, 16)), -- 15195 / 0x3b5b
    3170 => std_logic_vector(to_unsigned(12136, 16)), -- 12136 / 0x2f68 -- last item of row
    3171 => std_logic_vector(to_unsigned(   69, 16)), --    69 / 0x0045
    3172 => std_logic_vector(to_unsigned( 7758, 16)), --  7758 / 0x1e4e
    3173 => std_logic_vector(to_unsigned(22808, 16)), -- 22808 / 0x5918 -- last item of row
    3174 => std_logic_vector(to_unsigned(   70, 16)), --    70 / 0x0046
    3175 => std_logic_vector(to_unsigned( 3564, 16)), --  3564 / 0x0dec
    3176 => std_logic_vector(to_unsigned( 2925, 16)), --  2925 / 0x0b6d -- last item of row
    3177 => std_logic_vector(to_unsigned(   71, 16)), --    71 / 0x0047
    3178 => std_logic_vector(to_unsigned( 3434, 16)), --  3434 / 0x0d6a
    3179 => std_logic_vector(to_unsigned( 7769, 16)), --  7769 / 0x1e59 -- last item of row
    -- Table for fecframe_normal, C4_5
    3180 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3181 => std_logic_vector(to_unsigned(  149, 16)), --   149 / 0x0095
    3182 => std_logic_vector(to_unsigned(11212, 16)), -- 11212 / 0x2bcc
    3183 => std_logic_vector(to_unsigned( 5575, 16)), --  5575 / 0x15c7
    3184 => std_logic_vector(to_unsigned( 6360, 16)), --  6360 / 0x18d8
    3185 => std_logic_vector(to_unsigned(12559, 16)), -- 12559 / 0x310f
    3186 => std_logic_vector(to_unsigned( 8108, 16)), --  8108 / 0x1fac
    3187 => std_logic_vector(to_unsigned( 8505, 16)), --  8505 / 0x2139
    3188 => std_logic_vector(to_unsigned(  408, 16)), --   408 / 0x0198
    3189 => std_logic_vector(to_unsigned(10026, 16)), -- 10026 / 0x272a
    3190 => std_logic_vector(to_unsigned(12828, 16)), -- 12828 / 0x321c -- last item of row
    3191 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    3192 => std_logic_vector(to_unsigned( 5237, 16)), --  5237 / 0x1475
    3193 => std_logic_vector(to_unsigned(  490, 16)), --   490 / 0x01ea
    3194 => std_logic_vector(to_unsigned(10677, 16)), -- 10677 / 0x29b5
    3195 => std_logic_vector(to_unsigned( 4998, 16)), --  4998 / 0x1386
    3196 => std_logic_vector(to_unsigned( 3869, 16)), --  3869 / 0x0f1d
    3197 => std_logic_vector(to_unsigned( 3734, 16)), --  3734 / 0x0e96
    3198 => std_logic_vector(to_unsigned( 3092, 16)), --  3092 / 0x0c14
    3199 => std_logic_vector(to_unsigned( 3509, 16)), --  3509 / 0x0db5
    3200 => std_logic_vector(to_unsigned( 7703, 16)), --  7703 / 0x1e17
    3201 => std_logic_vector(to_unsigned(10305, 16)), -- 10305 / 0x2841 -- last item of row
    3202 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    3203 => std_logic_vector(to_unsigned( 8742, 16)), --  8742 / 0x2226
    3204 => std_logic_vector(to_unsigned( 5553, 16)), --  5553 / 0x15b1
    3205 => std_logic_vector(to_unsigned( 2820, 16)), --  2820 / 0x0b04
    3206 => std_logic_vector(to_unsigned( 7085, 16)), --  7085 / 0x1bad
    3207 => std_logic_vector(to_unsigned(12116, 16)), -- 12116 / 0x2f54
    3208 => std_logic_vector(to_unsigned(10485, 16)), -- 10485 / 0x28f5
    3209 => std_logic_vector(to_unsigned(  564, 16)), --   564 / 0x0234
    3210 => std_logic_vector(to_unsigned( 7795, 16)), --  7795 / 0x1e73
    3211 => std_logic_vector(to_unsigned( 2972, 16)), --  2972 / 0x0b9c
    3212 => std_logic_vector(to_unsigned( 2157, 16)), --  2157 / 0x086d -- last item of row
    3213 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    3214 => std_logic_vector(to_unsigned( 2699, 16)), --  2699 / 0x0a8b
    3215 => std_logic_vector(to_unsigned( 4304, 16)), --  4304 / 0x10d0
    3216 => std_logic_vector(to_unsigned( 8350, 16)), --  8350 / 0x209e
    3217 => std_logic_vector(to_unsigned(  712, 16)), --   712 / 0x02c8
    3218 => std_logic_vector(to_unsigned( 2841, 16)), --  2841 / 0x0b19
    3219 => std_logic_vector(to_unsigned( 3250, 16)), --  3250 / 0x0cb2
    3220 => std_logic_vector(to_unsigned( 4731, 16)), --  4731 / 0x127b
    3221 => std_logic_vector(to_unsigned(10105, 16)), -- 10105 / 0x2779
    3222 => std_logic_vector(to_unsigned(  517, 16)), --   517 / 0x0205
    3223 => std_logic_vector(to_unsigned( 7516, 16)), --  7516 / 0x1d5c -- last item of row
    3224 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    3225 => std_logic_vector(to_unsigned(12067, 16)), -- 12067 / 0x2f23
    3226 => std_logic_vector(to_unsigned( 1351, 16)), --  1351 / 0x0547
    3227 => std_logic_vector(to_unsigned(11992, 16)), -- 11992 / 0x2ed8
    3228 => std_logic_vector(to_unsigned(12191, 16)), -- 12191 / 0x2f9f
    3229 => std_logic_vector(to_unsigned(11267, 16)), -- 11267 / 0x2c03
    3230 => std_logic_vector(to_unsigned( 5161, 16)), --  5161 / 0x1429
    3231 => std_logic_vector(to_unsigned(  537, 16)), --   537 / 0x0219
    3232 => std_logic_vector(to_unsigned( 6166, 16)), --  6166 / 0x1816
    3233 => std_logic_vector(to_unsigned( 4246, 16)), --  4246 / 0x1096
    3234 => std_logic_vector(to_unsigned( 2363, 16)), --  2363 / 0x093b -- last item of row
    3235 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    3236 => std_logic_vector(to_unsigned( 6828, 16)), --  6828 / 0x1aac
    3237 => std_logic_vector(to_unsigned( 7107, 16)), --  7107 / 0x1bc3
    3238 => std_logic_vector(to_unsigned( 2127, 16)), --  2127 / 0x084f
    3239 => std_logic_vector(to_unsigned( 3724, 16)), --  3724 / 0x0e8c
    3240 => std_logic_vector(to_unsigned( 5743, 16)), --  5743 / 0x166f
    3241 => std_logic_vector(to_unsigned(11040, 16)), -- 11040 / 0x2b20
    3242 => std_logic_vector(to_unsigned(10756, 16)), -- 10756 / 0x2a04
    3243 => std_logic_vector(to_unsigned( 4073, 16)), --  4073 / 0x0fe9
    3244 => std_logic_vector(to_unsigned( 1011, 16)), --  1011 / 0x03f3
    3245 => std_logic_vector(to_unsigned( 3422, 16)), --  3422 / 0x0d5e -- last item of row
    3246 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    3247 => std_logic_vector(to_unsigned(11259, 16)), -- 11259 / 0x2bfb
    3248 => std_logic_vector(to_unsigned( 1216, 16)), --  1216 / 0x04c0
    3249 => std_logic_vector(to_unsigned( 9526, 16)), --  9526 / 0x2536
    3250 => std_logic_vector(to_unsigned( 1466, 16)), --  1466 / 0x05ba
    3251 => std_logic_vector(to_unsigned(10816, 16)), -- 10816 / 0x2a40
    3252 => std_logic_vector(to_unsigned(  940, 16)), --   940 / 0x03ac
    3253 => std_logic_vector(to_unsigned( 3744, 16)), --  3744 / 0x0ea0
    3254 => std_logic_vector(to_unsigned( 2815, 16)), --  2815 / 0x0aff
    3255 => std_logic_vector(to_unsigned(11506, 16)), -- 11506 / 0x2cf2
    3256 => std_logic_vector(to_unsigned(11573, 16)), -- 11573 / 0x2d35 -- last item of row
    3257 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    3258 => std_logic_vector(to_unsigned( 4549, 16)), --  4549 / 0x11c5
    3259 => std_logic_vector(to_unsigned(11507, 16)), -- 11507 / 0x2cf3
    3260 => std_logic_vector(to_unsigned( 1118, 16)), --  1118 / 0x045e
    3261 => std_logic_vector(to_unsigned( 1274, 16)), --  1274 / 0x04fa
    3262 => std_logic_vector(to_unsigned(11751, 16)), -- 11751 / 0x2de7
    3263 => std_logic_vector(to_unsigned( 5207, 16)), --  5207 / 0x1457
    3264 => std_logic_vector(to_unsigned( 7854, 16)), --  7854 / 0x1eae
    3265 => std_logic_vector(to_unsigned(12803, 16)), -- 12803 / 0x3203
    3266 => std_logic_vector(to_unsigned( 4047, 16)), --  4047 / 0x0fcf
    3267 => std_logic_vector(to_unsigned( 6484, 16)), --  6484 / 0x1954 -- last item of row
    3268 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    3269 => std_logic_vector(to_unsigned( 8430, 16)), --  8430 / 0x20ee
    3270 => std_logic_vector(to_unsigned( 4115, 16)), --  4115 / 0x1013
    3271 => std_logic_vector(to_unsigned( 9440, 16)), --  9440 / 0x24e0
    3272 => std_logic_vector(to_unsigned(  413, 16)), --   413 / 0x019d
    3273 => std_logic_vector(to_unsigned( 4455, 16)), --  4455 / 0x1167
    3274 => std_logic_vector(to_unsigned( 2262, 16)), --  2262 / 0x08d6
    3275 => std_logic_vector(to_unsigned( 7915, 16)), --  7915 / 0x1eeb
    3276 => std_logic_vector(to_unsigned(12402, 16)), -- 12402 / 0x3072
    3277 => std_logic_vector(to_unsigned( 8579, 16)), --  8579 / 0x2183
    3278 => std_logic_vector(to_unsigned( 7052, 16)), --  7052 / 0x1b8c -- last item of row
    3279 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    3280 => std_logic_vector(to_unsigned( 3885, 16)), --  3885 / 0x0f2d
    3281 => std_logic_vector(to_unsigned( 9126, 16)), --  9126 / 0x23a6
    3282 => std_logic_vector(to_unsigned( 5665, 16)), --  5665 / 0x1621
    3283 => std_logic_vector(to_unsigned( 4505, 16)), --  4505 / 0x1199
    3284 => std_logic_vector(to_unsigned( 2343, 16)), --  2343 / 0x0927
    3285 => std_logic_vector(to_unsigned(  253, 16)), --   253 / 0x00fd
    3286 => std_logic_vector(to_unsigned( 4707, 16)), --  4707 / 0x1263
    3287 => std_logic_vector(to_unsigned( 3742, 16)), --  3742 / 0x0e9e
    3288 => std_logic_vector(to_unsigned( 4166, 16)), --  4166 / 0x1046
    3289 => std_logic_vector(to_unsigned( 1556, 16)), --  1556 / 0x0614 -- last item of row
    3290 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    3291 => std_logic_vector(to_unsigned( 1704, 16)), --  1704 / 0x06a8
    3292 => std_logic_vector(to_unsigned( 8936, 16)), --  8936 / 0x22e8
    3293 => std_logic_vector(to_unsigned( 6775, 16)), --  6775 / 0x1a77
    3294 => std_logic_vector(to_unsigned( 8639, 16)), --  8639 / 0x21bf
    3295 => std_logic_vector(to_unsigned( 8179, 16)), --  8179 / 0x1ff3
    3296 => std_logic_vector(to_unsigned( 7954, 16)), --  7954 / 0x1f12
    3297 => std_logic_vector(to_unsigned( 8234, 16)), --  8234 / 0x202a
    3298 => std_logic_vector(to_unsigned( 7850, 16)), --  7850 / 0x1eaa
    3299 => std_logic_vector(to_unsigned( 8883, 16)), --  8883 / 0x22b3
    3300 => std_logic_vector(to_unsigned( 8713, 16)), --  8713 / 0x2209 -- last item of row
    3301 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    3302 => std_logic_vector(to_unsigned(11716, 16)), -- 11716 / 0x2dc4
    3303 => std_logic_vector(to_unsigned( 4344, 16)), --  4344 / 0x10f8
    3304 => std_logic_vector(to_unsigned( 9087, 16)), --  9087 / 0x237f
    3305 => std_logic_vector(to_unsigned(11264, 16)), -- 11264 / 0x2c00
    3306 => std_logic_vector(to_unsigned( 2274, 16)), --  2274 / 0x08e2
    3307 => std_logic_vector(to_unsigned( 8832, 16)), --  8832 / 0x2280
    3308 => std_logic_vector(to_unsigned( 9147, 16)), --  9147 / 0x23bb
    3309 => std_logic_vector(to_unsigned(11930, 16)), -- 11930 / 0x2e9a
    3310 => std_logic_vector(to_unsigned( 6054, 16)), --  6054 / 0x17a6
    3311 => std_logic_vector(to_unsigned( 5455, 16)), --  5455 / 0x154f -- last item of row
    3312 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3313 => std_logic_vector(to_unsigned( 7323, 16)), --  7323 / 0x1c9b
    3314 => std_logic_vector(to_unsigned( 3970, 16)), --  3970 / 0x0f82
    3315 => std_logic_vector(to_unsigned(10329, 16)), -- 10329 / 0x2859
    3316 => std_logic_vector(to_unsigned( 2170, 16)), --  2170 / 0x087a
    3317 => std_logic_vector(to_unsigned( 8262, 16)), --  8262 / 0x2046
    3318 => std_logic_vector(to_unsigned( 3854, 16)), --  3854 / 0x0f0e
    3319 => std_logic_vector(to_unsigned( 2087, 16)), --  2087 / 0x0827
    3320 => std_logic_vector(to_unsigned(12899, 16)), -- 12899 / 0x3263
    3321 => std_logic_vector(to_unsigned( 9497, 16)), --  9497 / 0x2519
    3322 => std_logic_vector(to_unsigned(11700, 16)), -- 11700 / 0x2db4 -- last item of row
    3323 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3324 => std_logic_vector(to_unsigned( 4418, 16)), --  4418 / 0x1142
    3325 => std_logic_vector(to_unsigned( 1467, 16)), --  1467 / 0x05bb
    3326 => std_logic_vector(to_unsigned( 2490, 16)), --  2490 / 0x09ba
    3327 => std_logic_vector(to_unsigned( 5841, 16)), --  5841 / 0x16d1
    3328 => std_logic_vector(to_unsigned(  817, 16)), --   817 / 0x0331
    3329 => std_logic_vector(to_unsigned(11453, 16)), -- 11453 / 0x2cbd
    3330 => std_logic_vector(to_unsigned(  533, 16)), --   533 / 0x0215
    3331 => std_logic_vector(to_unsigned(11217, 16)), -- 11217 / 0x2bd1
    3332 => std_logic_vector(to_unsigned(11962, 16)), -- 11962 / 0x2eba
    3333 => std_logic_vector(to_unsigned( 5251, 16)), --  5251 / 0x1483 -- last item of row
    3334 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3335 => std_logic_vector(to_unsigned( 1541, 16)), --  1541 / 0x0605
    3336 => std_logic_vector(to_unsigned( 4525, 16)), --  4525 / 0x11ad
    3337 => std_logic_vector(to_unsigned( 7976, 16)), --  7976 / 0x1f28
    3338 => std_logic_vector(to_unsigned( 3457, 16)), --  3457 / 0x0d81
    3339 => std_logic_vector(to_unsigned( 9536, 16)), --  9536 / 0x2540
    3340 => std_logic_vector(to_unsigned( 7725, 16)), --  7725 / 0x1e2d
    3341 => std_logic_vector(to_unsigned( 3788, 16)), --  3788 / 0x0ecc
    3342 => std_logic_vector(to_unsigned( 2982, 16)), --  2982 / 0x0ba6
    3343 => std_logic_vector(to_unsigned( 6307, 16)), --  6307 / 0x18a3
    3344 => std_logic_vector(to_unsigned( 5997, 16)), --  5997 / 0x176d -- last item of row
    3345 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3346 => std_logic_vector(to_unsigned(11484, 16)), -- 11484 / 0x2cdc
    3347 => std_logic_vector(to_unsigned( 2739, 16)), --  2739 / 0x0ab3
    3348 => std_logic_vector(to_unsigned( 4023, 16)), --  4023 / 0x0fb7
    3349 => std_logic_vector(to_unsigned(12107, 16)), -- 12107 / 0x2f4b
    3350 => std_logic_vector(to_unsigned( 6516, 16)), --  6516 / 0x1974
    3351 => std_logic_vector(to_unsigned(  551, 16)), --   551 / 0x0227
    3352 => std_logic_vector(to_unsigned( 2572, 16)), --  2572 / 0x0a0c
    3353 => std_logic_vector(to_unsigned( 6628, 16)), --  6628 / 0x19e4
    3354 => std_logic_vector(to_unsigned( 8150, 16)), --  8150 / 0x1fd6
    3355 => std_logic_vector(to_unsigned( 9852, 16)), --  9852 / 0x267c -- last item of row
    3356 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3357 => std_logic_vector(to_unsigned( 6070, 16)), --  6070 / 0x17b6
    3358 => std_logic_vector(to_unsigned( 1761, 16)), --  1761 / 0x06e1
    3359 => std_logic_vector(to_unsigned( 4627, 16)), --  4627 / 0x1213
    3360 => std_logic_vector(to_unsigned( 6534, 16)), --  6534 / 0x1986
    3361 => std_logic_vector(to_unsigned( 7913, 16)), --  7913 / 0x1ee9
    3362 => std_logic_vector(to_unsigned( 3730, 16)), --  3730 / 0x0e92
    3363 => std_logic_vector(to_unsigned(11866, 16)), -- 11866 / 0x2e5a
    3364 => std_logic_vector(to_unsigned( 1813, 16)), --  1813 / 0x0715
    3365 => std_logic_vector(to_unsigned(12306, 16)), -- 12306 / 0x3012
    3366 => std_logic_vector(to_unsigned( 8249, 16)), --  8249 / 0x2039 -- last item of row
    3367 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3368 => std_logic_vector(to_unsigned(12441, 16)), -- 12441 / 0x3099
    3369 => std_logic_vector(to_unsigned( 5489, 16)), --  5489 / 0x1571
    3370 => std_logic_vector(to_unsigned( 8748, 16)), --  8748 / 0x222c
    3371 => std_logic_vector(to_unsigned( 7837, 16)), --  7837 / 0x1e9d
    3372 => std_logic_vector(to_unsigned( 7660, 16)), --  7660 / 0x1dec
    3373 => std_logic_vector(to_unsigned( 2102, 16)), --  2102 / 0x0836
    3374 => std_logic_vector(to_unsigned(11341, 16)), -- 11341 / 0x2c4d
    3375 => std_logic_vector(to_unsigned( 2936, 16)), --  2936 / 0x0b78
    3376 => std_logic_vector(to_unsigned( 6712, 16)), --  6712 / 0x1a38
    3377 => std_logic_vector(to_unsigned(11977, 16)), -- 11977 / 0x2ec9 -- last item of row
    3378 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3379 => std_logic_vector(to_unsigned(10155, 16)), -- 10155 / 0x27ab
    3380 => std_logic_vector(to_unsigned( 4210, 16)), --  4210 / 0x1072 -- last item of row
    3381 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3382 => std_logic_vector(to_unsigned( 1010, 16)), --  1010 / 0x03f2
    3383 => std_logic_vector(to_unsigned(10483, 16)), -- 10483 / 0x28f3 -- last item of row
    3384 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3385 => std_logic_vector(to_unsigned( 8900, 16)), --  8900 / 0x22c4
    3386 => std_logic_vector(to_unsigned(10250, 16)), -- 10250 / 0x280a -- last item of row
    3387 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3388 => std_logic_vector(to_unsigned(10243, 16)), -- 10243 / 0x2803
    3389 => std_logic_vector(to_unsigned(12278, 16)), -- 12278 / 0x2ff6 -- last item of row
    3390 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3391 => std_logic_vector(to_unsigned( 7070, 16)), --  7070 / 0x1b9e
    3392 => std_logic_vector(to_unsigned( 4397, 16)), --  4397 / 0x112d -- last item of row
    3393 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3394 => std_logic_vector(to_unsigned(12271, 16)), -- 12271 / 0x2fef
    3395 => std_logic_vector(to_unsigned( 3887, 16)), --  3887 / 0x0f2f -- last item of row
    3396 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3397 => std_logic_vector(to_unsigned(11980, 16)), -- 11980 / 0x2ecc
    3398 => std_logic_vector(to_unsigned( 6836, 16)), --  6836 / 0x1ab4 -- last item of row
    3399 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3400 => std_logic_vector(to_unsigned( 9514, 16)), --  9514 / 0x252a
    3401 => std_logic_vector(to_unsigned( 4356, 16)), --  4356 / 0x1104 -- last item of row
    3402 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3403 => std_logic_vector(to_unsigned( 7137, 16)), --  7137 / 0x1be1
    3404 => std_logic_vector(to_unsigned(10281, 16)), -- 10281 / 0x2829 -- last item of row
    3405 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3406 => std_logic_vector(to_unsigned(11881, 16)), -- 11881 / 0x2e69
    3407 => std_logic_vector(to_unsigned( 2526, 16)), --  2526 / 0x09de -- last item of row
    3408 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3409 => std_logic_vector(to_unsigned( 1969, 16)), --  1969 / 0x07b1
    3410 => std_logic_vector(to_unsigned(11477, 16)), -- 11477 / 0x2cd5 -- last item of row
    3411 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3412 => std_logic_vector(to_unsigned( 3044, 16)), --  3044 / 0x0be4
    3413 => std_logic_vector(to_unsigned(10921, 16)), -- 10921 / 0x2aa9 -- last item of row
    3414 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    3415 => std_logic_vector(to_unsigned( 2236, 16)), --  2236 / 0x08bc
    3416 => std_logic_vector(to_unsigned( 8724, 16)), --  8724 / 0x2214 -- last item of row
    3417 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    3418 => std_logic_vector(to_unsigned( 9104, 16)), --  9104 / 0x2390
    3419 => std_logic_vector(to_unsigned( 6340, 16)), --  6340 / 0x18c4 -- last item of row
    3420 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    3421 => std_logic_vector(to_unsigned( 7342, 16)), --  7342 / 0x1cae
    3422 => std_logic_vector(to_unsigned( 8582, 16)), --  8582 / 0x2186 -- last item of row
    3423 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    3424 => std_logic_vector(to_unsigned(11675, 16)), -- 11675 / 0x2d9b
    3425 => std_logic_vector(to_unsigned(10405, 16)), -- 10405 / 0x28a5 -- last item of row
    3426 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    3427 => std_logic_vector(to_unsigned( 6467, 16)), --  6467 / 0x1943
    3428 => std_logic_vector(to_unsigned(12775, 16)), -- 12775 / 0x31e7 -- last item of row
    3429 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    3430 => std_logic_vector(to_unsigned( 3186, 16)), --  3186 / 0x0c72
    3431 => std_logic_vector(to_unsigned(12198, 16)), -- 12198 / 0x2fa6 -- last item of row
    3432 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3433 => std_logic_vector(to_unsigned( 9621, 16)), --  9621 / 0x2595
    3434 => std_logic_vector(to_unsigned(11445, 16)), -- 11445 / 0x2cb5 -- last item of row
    3435 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    3436 => std_logic_vector(to_unsigned( 7486, 16)), --  7486 / 0x1d3e
    3437 => std_logic_vector(to_unsigned( 5611, 16)), --  5611 / 0x15eb -- last item of row
    3438 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    3439 => std_logic_vector(to_unsigned( 4319, 16)), --  4319 / 0x10df
    3440 => std_logic_vector(to_unsigned( 4879, 16)), --  4879 / 0x130f -- last item of row
    3441 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    3442 => std_logic_vector(to_unsigned( 2196, 16)), --  2196 / 0x0894
    3443 => std_logic_vector(to_unsigned(  344, 16)), --   344 / 0x0158 -- last item of row
    3444 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    3445 => std_logic_vector(to_unsigned( 7527, 16)), --  7527 / 0x1d67
    3446 => std_logic_vector(to_unsigned( 6650, 16)), --  6650 / 0x19fa -- last item of row
    3447 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    3448 => std_logic_vector(to_unsigned(10693, 16)), -- 10693 / 0x29c5
    3449 => std_logic_vector(to_unsigned( 2440, 16)), --  2440 / 0x0988 -- last item of row
    3450 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    3451 => std_logic_vector(to_unsigned( 6755, 16)), --  6755 / 0x1a63
    3452 => std_logic_vector(to_unsigned( 2706, 16)), --  2706 / 0x0a92 -- last item of row
    3453 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    3454 => std_logic_vector(to_unsigned( 5144, 16)), --  5144 / 0x1418
    3455 => std_logic_vector(to_unsigned( 5998, 16)), --  5998 / 0x176e -- last item of row
    3456 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    3457 => std_logic_vector(to_unsigned(11043, 16)), -- 11043 / 0x2b23
    3458 => std_logic_vector(to_unsigned( 8033, 16)), --  8033 / 0x1f61 -- last item of row
    3459 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    3460 => std_logic_vector(to_unsigned( 4846, 16)), --  4846 / 0x12ee
    3461 => std_logic_vector(to_unsigned( 4435, 16)), --  4435 / 0x1153 -- last item of row
    3462 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    3463 => std_logic_vector(to_unsigned( 4157, 16)), --  4157 / 0x103d
    3464 => std_logic_vector(to_unsigned( 9228, 16)), --  9228 / 0x240c -- last item of row
    3465 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    3466 => std_logic_vector(to_unsigned(12270, 16)), -- 12270 / 0x2fee
    3467 => std_logic_vector(to_unsigned( 6562, 16)), --  6562 / 0x19a2 -- last item of row
    3468 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3469 => std_logic_vector(to_unsigned(11954, 16)), -- 11954 / 0x2eb2
    3470 => std_logic_vector(to_unsigned( 7592, 16)), --  7592 / 0x1da8 -- last item of row
    3471 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3472 => std_logic_vector(to_unsigned( 7420, 16)), --  7420 / 0x1cfc
    3473 => std_logic_vector(to_unsigned( 2592, 16)), --  2592 / 0x0a20 -- last item of row
    3474 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3475 => std_logic_vector(to_unsigned( 8810, 16)), --  8810 / 0x226a
    3476 => std_logic_vector(to_unsigned( 9636, 16)), --  9636 / 0x25a4 -- last item of row
    3477 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3478 => std_logic_vector(to_unsigned(  689, 16)), --   689 / 0x02b1
    3479 => std_logic_vector(to_unsigned( 5430, 16)), --  5430 / 0x1536 -- last item of row
    3480 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3481 => std_logic_vector(to_unsigned(  920, 16)), --   920 / 0x0398
    3482 => std_logic_vector(to_unsigned( 1304, 16)), --  1304 / 0x0518 -- last item of row
    3483 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3484 => std_logic_vector(to_unsigned( 1253, 16)), --  1253 / 0x04e5
    3485 => std_logic_vector(to_unsigned(11934, 16)), -- 11934 / 0x2e9e -- last item of row
    3486 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3487 => std_logic_vector(to_unsigned( 9559, 16)), --  9559 / 0x2557
    3488 => std_logic_vector(to_unsigned( 6016, 16)), --  6016 / 0x1780 -- last item of row
    3489 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3490 => std_logic_vector(to_unsigned(  312, 16)), --   312 / 0x0138
    3491 => std_logic_vector(to_unsigned( 7589, 16)), --  7589 / 0x1da5 -- last item of row
    3492 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3493 => std_logic_vector(to_unsigned( 4439, 16)), --  4439 / 0x1157
    3494 => std_logic_vector(to_unsigned( 4197, 16)), --  4197 / 0x1065 -- last item of row
    3495 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3496 => std_logic_vector(to_unsigned( 4002, 16)), --  4002 / 0x0fa2
    3497 => std_logic_vector(to_unsigned( 9555, 16)), --  9555 / 0x2553 -- last item of row
    3498 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3499 => std_logic_vector(to_unsigned(12232, 16)), -- 12232 / 0x2fc8
    3500 => std_logic_vector(to_unsigned( 7779, 16)), --  7779 / 0x1e63 -- last item of row
    3501 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3502 => std_logic_vector(to_unsigned( 1494, 16)), --  1494 / 0x05d6
    3503 => std_logic_vector(to_unsigned( 8782, 16)), --  8782 / 0x224e -- last item of row
    3504 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3505 => std_logic_vector(to_unsigned(10749, 16)), -- 10749 / 0x29fd
    3506 => std_logic_vector(to_unsigned( 3969, 16)), --  3969 / 0x0f81 -- last item of row
    3507 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3508 => std_logic_vector(to_unsigned( 4368, 16)), --  4368 / 0x1110
    3509 => std_logic_vector(to_unsigned( 3479, 16)), --  3479 / 0x0d97 -- last item of row
    3510 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3511 => std_logic_vector(to_unsigned( 6316, 16)), --  6316 / 0x18ac
    3512 => std_logic_vector(to_unsigned( 5342, 16)), --  5342 / 0x14de -- last item of row
    3513 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3514 => std_logic_vector(to_unsigned( 2455, 16)), --  2455 / 0x0997
    3515 => std_logic_vector(to_unsigned( 3493, 16)), --  3493 / 0x0da5 -- last item of row
    3516 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3517 => std_logic_vector(to_unsigned(12157, 16)), -- 12157 / 0x2f7d
    3518 => std_logic_vector(to_unsigned( 7405, 16)), --  7405 / 0x1ced -- last item of row
    3519 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3520 => std_logic_vector(to_unsigned( 6598, 16)), --  6598 / 0x19c6
    3521 => std_logic_vector(to_unsigned(11495, 16)), -- 11495 / 0x2ce7 -- last item of row
    3522 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    3523 => std_logic_vector(to_unsigned(11805, 16)), -- 11805 / 0x2e1d
    3524 => std_logic_vector(to_unsigned( 4455, 16)), --  4455 / 0x1167 -- last item of row
    3525 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    3526 => std_logic_vector(to_unsigned( 9625, 16)), --  9625 / 0x2599
    3527 => std_logic_vector(to_unsigned( 2090, 16)), --  2090 / 0x082a -- last item of row
    3528 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    3529 => std_logic_vector(to_unsigned( 4731, 16)), --  4731 / 0x127b
    3530 => std_logic_vector(to_unsigned( 2321, 16)), --  2321 / 0x0911 -- last item of row
    3531 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    3532 => std_logic_vector(to_unsigned( 3578, 16)), --  3578 / 0x0dfa
    3533 => std_logic_vector(to_unsigned( 2608, 16)), --  2608 / 0x0a30 -- last item of row
    3534 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    3535 => std_logic_vector(to_unsigned( 8504, 16)), --  8504 / 0x2138
    3536 => std_logic_vector(to_unsigned( 1849, 16)), --  1849 / 0x0739 -- last item of row
    3537 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    3538 => std_logic_vector(to_unsigned( 4027, 16)), --  4027 / 0x0fbb
    3539 => std_logic_vector(to_unsigned( 1151, 16)), --  1151 / 0x047f -- last item of row
    3540 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3541 => std_logic_vector(to_unsigned( 5647, 16)), --  5647 / 0x160f
    3542 => std_logic_vector(to_unsigned( 4935, 16)), --  4935 / 0x1347 -- last item of row
    3543 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    3544 => std_logic_vector(to_unsigned( 4219, 16)), --  4219 / 0x107b
    3545 => std_logic_vector(to_unsigned( 1870, 16)), --  1870 / 0x074e -- last item of row
    3546 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    3547 => std_logic_vector(to_unsigned(10968, 16)), -- 10968 / 0x2ad8
    3548 => std_logic_vector(to_unsigned( 8054, 16)), --  8054 / 0x1f76 -- last item of row
    3549 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    3550 => std_logic_vector(to_unsigned( 6970, 16)), --  6970 / 0x1b3a
    3551 => std_logic_vector(to_unsigned( 5447, 16)), --  5447 / 0x1547 -- last item of row
    3552 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    3553 => std_logic_vector(to_unsigned( 3217, 16)), --  3217 / 0x0c91
    3554 => std_logic_vector(to_unsigned( 5638, 16)), --  5638 / 0x1606 -- last item of row
    3555 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    3556 => std_logic_vector(to_unsigned( 8972, 16)), --  8972 / 0x230c
    3557 => std_logic_vector(to_unsigned(  669, 16)), --   669 / 0x029d -- last item of row
    3558 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    3559 => std_logic_vector(to_unsigned( 5618, 16)), --  5618 / 0x15f2
    3560 => std_logic_vector(to_unsigned(12472, 16)), -- 12472 / 0x30b8 -- last item of row
    3561 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    3562 => std_logic_vector(to_unsigned( 1457, 16)), --  1457 / 0x05b1
    3563 => std_logic_vector(to_unsigned( 1280, 16)), --  1280 / 0x0500 -- last item of row
    3564 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    3565 => std_logic_vector(to_unsigned( 8868, 16)), --  8868 / 0x22a4
    3566 => std_logic_vector(to_unsigned( 3883, 16)), --  3883 / 0x0f2b -- last item of row
    3567 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    3568 => std_logic_vector(to_unsigned( 8866, 16)), --  8866 / 0x22a2
    3569 => std_logic_vector(to_unsigned( 1224, 16)), --  1224 / 0x04c8 -- last item of row
    3570 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    3571 => std_logic_vector(to_unsigned( 8371, 16)), --  8371 / 0x20b3
    3572 => std_logic_vector(to_unsigned( 5972, 16)), --  5972 / 0x1754 -- last item of row
    3573 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    3574 => std_logic_vector(to_unsigned(  266, 16)), --   266 / 0x010a
    3575 => std_logic_vector(to_unsigned( 4405, 16)), --  4405 / 0x1135 -- last item of row
    3576 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3577 => std_logic_vector(to_unsigned( 3706, 16)), --  3706 / 0x0e7a
    3578 => std_logic_vector(to_unsigned( 3244, 16)), --  3244 / 0x0cac -- last item of row
    3579 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3580 => std_logic_vector(to_unsigned( 6039, 16)), --  6039 / 0x1797
    3581 => std_logic_vector(to_unsigned( 5844, 16)), --  5844 / 0x16d4 -- last item of row
    3582 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3583 => std_logic_vector(to_unsigned( 7200, 16)), --  7200 / 0x1c20
    3584 => std_logic_vector(to_unsigned( 3283, 16)), --  3283 / 0x0cd3 -- last item of row
    3585 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3586 => std_logic_vector(to_unsigned( 1502, 16)), --  1502 / 0x05de
    3587 => std_logic_vector(to_unsigned(11282, 16)), -- 11282 / 0x2c12 -- last item of row
    3588 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3589 => std_logic_vector(to_unsigned(12318, 16)), -- 12318 / 0x301e
    3590 => std_logic_vector(to_unsigned( 2202, 16)), --  2202 / 0x089a -- last item of row
    3591 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3592 => std_logic_vector(to_unsigned( 4523, 16)), --  4523 / 0x11ab
    3593 => std_logic_vector(to_unsigned(  965, 16)), --   965 / 0x03c5 -- last item of row
    3594 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3595 => std_logic_vector(to_unsigned( 9587, 16)), --  9587 / 0x2573
    3596 => std_logic_vector(to_unsigned( 7011, 16)), --  7011 / 0x1b63 -- last item of row
    3597 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3598 => std_logic_vector(to_unsigned( 2552, 16)), --  2552 / 0x09f8
    3599 => std_logic_vector(to_unsigned( 2051, 16)), --  2051 / 0x0803 -- last item of row
    3600 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3601 => std_logic_vector(to_unsigned(12045, 16)), -- 12045 / 0x2f0d
    3602 => std_logic_vector(to_unsigned(10306, 16)), -- 10306 / 0x2842 -- last item of row
    3603 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3604 => std_logic_vector(to_unsigned(11070, 16)), -- 11070 / 0x2b3e
    3605 => std_logic_vector(to_unsigned( 5104, 16)), --  5104 / 0x13f0 -- last item of row
    3606 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3607 => std_logic_vector(to_unsigned( 6627, 16)), --  6627 / 0x19e3
    3608 => std_logic_vector(to_unsigned( 6906, 16)), --  6906 / 0x1afa -- last item of row
    3609 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3610 => std_logic_vector(to_unsigned( 9889, 16)), --  9889 / 0x26a1
    3611 => std_logic_vector(to_unsigned( 2121, 16)), --  2121 / 0x0849 -- last item of row
    3612 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3613 => std_logic_vector(to_unsigned(  829, 16)), --   829 / 0x033d
    3614 => std_logic_vector(to_unsigned( 9701, 16)), --  9701 / 0x25e5 -- last item of row
    3615 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3616 => std_logic_vector(to_unsigned( 2201, 16)), --  2201 / 0x0899
    3617 => std_logic_vector(to_unsigned( 1819, 16)), --  1819 / 0x071b -- last item of row
    3618 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3619 => std_logic_vector(to_unsigned( 6689, 16)), --  6689 / 0x1a21
    3620 => std_logic_vector(to_unsigned(12925, 16)), -- 12925 / 0x327d -- last item of row
    3621 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3622 => std_logic_vector(to_unsigned( 2139, 16)), --  2139 / 0x085b
    3623 => std_logic_vector(to_unsigned( 8757, 16)), --  8757 / 0x2235 -- last item of row
    3624 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3625 => std_logic_vector(to_unsigned(12004, 16)), -- 12004 / 0x2ee4
    3626 => std_logic_vector(to_unsigned( 5948, 16)), --  5948 / 0x173c -- last item of row
    3627 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3628 => std_logic_vector(to_unsigned( 8704, 16)), --  8704 / 0x2200
    3629 => std_logic_vector(to_unsigned( 3191, 16)), --  3191 / 0x0c77 -- last item of row
    3630 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    3631 => std_logic_vector(to_unsigned( 8171, 16)), --  8171 / 0x1feb
    3632 => std_logic_vector(to_unsigned(10933, 16)), -- 10933 / 0x2ab5 -- last item of row
    3633 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    3634 => std_logic_vector(to_unsigned( 6297, 16)), --  6297 / 0x1899
    3635 => std_logic_vector(to_unsigned( 7116, 16)), --  7116 / 0x1bcc -- last item of row
    3636 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    3637 => std_logic_vector(to_unsigned(  616, 16)), --   616 / 0x0268
    3638 => std_logic_vector(to_unsigned( 7146, 16)), --  7146 / 0x1bea -- last item of row
    3639 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    3640 => std_logic_vector(to_unsigned( 5142, 16)), --  5142 / 0x1416
    3641 => std_logic_vector(to_unsigned( 9761, 16)), --  9761 / 0x2621 -- last item of row
    3642 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    3643 => std_logic_vector(to_unsigned(10377, 16)), -- 10377 / 0x2889
    3644 => std_logic_vector(to_unsigned( 8138, 16)), --  8138 / 0x1fca -- last item of row
    3645 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    3646 => std_logic_vector(to_unsigned( 7616, 16)), --  7616 / 0x1dc0
    3647 => std_logic_vector(to_unsigned( 5811, 16)), --  5811 / 0x16b3 -- last item of row
    3648 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3649 => std_logic_vector(to_unsigned( 7285, 16)), --  7285 / 0x1c75
    3650 => std_logic_vector(to_unsigned( 9863, 16)), --  9863 / 0x2687 -- last item of row
    3651 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    3652 => std_logic_vector(to_unsigned( 7764, 16)), --  7764 / 0x1e54
    3653 => std_logic_vector(to_unsigned(10867, 16)), -- 10867 / 0x2a73 -- last item of row
    3654 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    3655 => std_logic_vector(to_unsigned(12343, 16)), -- 12343 / 0x3037
    3656 => std_logic_vector(to_unsigned( 9019, 16)), --  9019 / 0x233b -- last item of row
    3657 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    3658 => std_logic_vector(to_unsigned( 4414, 16)), --  4414 / 0x113e
    3659 => std_logic_vector(to_unsigned( 8331, 16)), --  8331 / 0x208b -- last item of row
    3660 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    3661 => std_logic_vector(to_unsigned( 3464, 16)), --  3464 / 0x0d88
    3662 => std_logic_vector(to_unsigned(  642, 16)), --   642 / 0x0282 -- last item of row
    3663 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    3664 => std_logic_vector(to_unsigned( 6960, 16)), --  6960 / 0x1b30
    3665 => std_logic_vector(to_unsigned( 2039, 16)), --  2039 / 0x07f7 -- last item of row
    3666 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    3667 => std_logic_vector(to_unsigned(  786, 16)), --   786 / 0x0312
    3668 => std_logic_vector(to_unsigned( 3021, 16)), --  3021 / 0x0bcd -- last item of row
    3669 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    3670 => std_logic_vector(to_unsigned(  710, 16)), --   710 / 0x02c6
    3671 => std_logic_vector(to_unsigned( 2086, 16)), --  2086 / 0x0826 -- last item of row
    3672 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    3673 => std_logic_vector(to_unsigned( 7423, 16)), --  7423 / 0x1cff
    3674 => std_logic_vector(to_unsigned( 5601, 16)), --  5601 / 0x15e1 -- last item of row
    3675 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    3676 => std_logic_vector(to_unsigned( 8120, 16)), --  8120 / 0x1fb8
    3677 => std_logic_vector(to_unsigned( 4885, 16)), --  4885 / 0x1315 -- last item of row
    3678 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    3679 => std_logic_vector(to_unsigned(12385, 16)), -- 12385 / 0x3061
    3680 => std_logic_vector(to_unsigned(11990, 16)), -- 11990 / 0x2ed6 -- last item of row
    3681 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    3682 => std_logic_vector(to_unsigned( 9739, 16)), --  9739 / 0x260b
    3683 => std_logic_vector(to_unsigned(10034, 16)), -- 10034 / 0x2732 -- last item of row
    3684 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3685 => std_logic_vector(to_unsigned(  424, 16)), --   424 / 0x01a8
    3686 => std_logic_vector(to_unsigned(10162, 16)), -- 10162 / 0x27b2 -- last item of row
    3687 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3688 => std_logic_vector(to_unsigned( 1347, 16)), --  1347 / 0x0543
    3689 => std_logic_vector(to_unsigned( 7597, 16)), --  7597 / 0x1dad -- last item of row
    3690 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3691 => std_logic_vector(to_unsigned( 1450, 16)), --  1450 / 0x05aa
    3692 => std_logic_vector(to_unsigned(  112, 16)), --   112 / 0x0070 -- last item of row
    3693 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3694 => std_logic_vector(to_unsigned( 7965, 16)), --  7965 / 0x1f1d
    3695 => std_logic_vector(to_unsigned( 8478, 16)), --  8478 / 0x211e -- last item of row
    3696 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3697 => std_logic_vector(to_unsigned( 8945, 16)), --  8945 / 0x22f1
    3698 => std_logic_vector(to_unsigned( 7397, 16)), --  7397 / 0x1ce5 -- last item of row
    3699 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3700 => std_logic_vector(to_unsigned( 6590, 16)), --  6590 / 0x19be
    3701 => std_logic_vector(to_unsigned( 8316, 16)), --  8316 / 0x207c -- last item of row
    3702 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3703 => std_logic_vector(to_unsigned( 6838, 16)), --  6838 / 0x1ab6
    3704 => std_logic_vector(to_unsigned( 9011, 16)), --  9011 / 0x2333 -- last item of row
    3705 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3706 => std_logic_vector(to_unsigned( 6174, 16)), --  6174 / 0x181e
    3707 => std_logic_vector(to_unsigned( 9410, 16)), --  9410 / 0x24c2 -- last item of row
    3708 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3709 => std_logic_vector(to_unsigned(  255, 16)), --   255 / 0x00ff
    3710 => std_logic_vector(to_unsigned(  113, 16)), --   113 / 0x0071 -- last item of row
    3711 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3712 => std_logic_vector(to_unsigned( 6197, 16)), --  6197 / 0x1835
    3713 => std_logic_vector(to_unsigned( 5835, 16)), --  5835 / 0x16cb -- last item of row
    3714 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3715 => std_logic_vector(to_unsigned(12902, 16)), -- 12902 / 0x3266
    3716 => std_logic_vector(to_unsigned( 3844, 16)), --  3844 / 0x0f04 -- last item of row
    3717 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3718 => std_logic_vector(to_unsigned( 4377, 16)), --  4377 / 0x1119
    3719 => std_logic_vector(to_unsigned( 3505, 16)), --  3505 / 0x0db1 -- last item of row
    3720 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3721 => std_logic_vector(to_unsigned( 5478, 16)), --  5478 / 0x1566
    3722 => std_logic_vector(to_unsigned( 8672, 16)), --  8672 / 0x21e0 -- last item of row
    3723 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3724 => std_logic_vector(to_unsigned( 4453, 16)), --  4453 / 0x1165
    3725 => std_logic_vector(to_unsigned( 2132, 16)), --  2132 / 0x0854 -- last item of row
    3726 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3727 => std_logic_vector(to_unsigned( 9724, 16)), --  9724 / 0x25fc
    3728 => std_logic_vector(to_unsigned( 1380, 16)), --  1380 / 0x0564 -- last item of row
    3729 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3730 => std_logic_vector(to_unsigned(12131, 16)), -- 12131 / 0x2f63
    3731 => std_logic_vector(to_unsigned(11526, 16)), -- 11526 / 0x2d06 -- last item of row
    3732 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3733 => std_logic_vector(to_unsigned(12323, 16)), -- 12323 / 0x3023
    3734 => std_logic_vector(to_unsigned( 9511, 16)), --  9511 / 0x2527 -- last item of row
    3735 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3736 => std_logic_vector(to_unsigned( 8231, 16)), --  8231 / 0x2027
    3737 => std_logic_vector(to_unsigned( 1752, 16)), --  1752 / 0x06d8 -- last item of row
    3738 => std_logic_vector(to_unsigned(   30, 16)), --    30 / 0x001e
    3739 => std_logic_vector(to_unsigned(  497, 16)), --   497 / 0x01f1
    3740 => std_logic_vector(to_unsigned( 9022, 16)), --  9022 / 0x233e -- last item of row
    3741 => std_logic_vector(to_unsigned(   31, 16)), --    31 / 0x001f
    3742 => std_logic_vector(to_unsigned( 9288, 16)), --  9288 / 0x2448
    3743 => std_logic_vector(to_unsigned( 3080, 16)), --  3080 / 0x0c08 -- last item of row
    3744 => std_logic_vector(to_unsigned(   32, 16)), --    32 / 0x0020
    3745 => std_logic_vector(to_unsigned( 2481, 16)), --  2481 / 0x09b1
    3746 => std_logic_vector(to_unsigned( 7515, 16)), --  7515 / 0x1d5b -- last item of row
    3747 => std_logic_vector(to_unsigned(   33, 16)), --    33 / 0x0021
    3748 => std_logic_vector(to_unsigned( 2696, 16)), --  2696 / 0x0a88
    3749 => std_logic_vector(to_unsigned(  268, 16)), --   268 / 0x010c -- last item of row
    3750 => std_logic_vector(to_unsigned(   34, 16)), --    34 / 0x0022
    3751 => std_logic_vector(to_unsigned( 4023, 16)), --  4023 / 0x0fb7
    3752 => std_logic_vector(to_unsigned(12341, 16)), -- 12341 / 0x3035 -- last item of row
    3753 => std_logic_vector(to_unsigned(   35, 16)), --    35 / 0x0023
    3754 => std_logic_vector(to_unsigned( 7108, 16)), --  7108 / 0x1bc4
    3755 => std_logic_vector(to_unsigned( 5553, 16)), --  5553 / 0x15b1 -- last item of row
    -- Table for fecframe_normal, C5_6
    3756 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3757 => std_logic_vector(to_unsigned( 4362, 16)), --  4362 / 0x110a
    3758 => std_logic_vector(to_unsigned(  416, 16)), --   416 / 0x01a0
    3759 => std_logic_vector(to_unsigned( 8909, 16)), --  8909 / 0x22cd
    3760 => std_logic_vector(to_unsigned( 4156, 16)), --  4156 / 0x103c
    3761 => std_logic_vector(to_unsigned( 3216, 16)), --  3216 / 0x0c90
    3762 => std_logic_vector(to_unsigned( 3112, 16)), --  3112 / 0x0c28
    3763 => std_logic_vector(to_unsigned( 2560, 16)), --  2560 / 0x0a00
    3764 => std_logic_vector(to_unsigned( 2912, 16)), --  2912 / 0x0b60
    3765 => std_logic_vector(to_unsigned( 6405, 16)), --  6405 / 0x1905
    3766 => std_logic_vector(to_unsigned( 8593, 16)), --  8593 / 0x2191
    3767 => std_logic_vector(to_unsigned( 4969, 16)), --  4969 / 0x1369
    3768 => std_logic_vector(to_unsigned( 6723, 16)), --  6723 / 0x1a43 -- last item of row
    3769 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    3770 => std_logic_vector(to_unsigned( 2479, 16)), --  2479 / 0x09af
    3771 => std_logic_vector(to_unsigned( 1786, 16)), --  1786 / 0x06fa
    3772 => std_logic_vector(to_unsigned( 8978, 16)), --  8978 / 0x2312
    3773 => std_logic_vector(to_unsigned( 3011, 16)), --  3011 / 0x0bc3
    3774 => std_logic_vector(to_unsigned( 4339, 16)), --  4339 / 0x10f3
    3775 => std_logic_vector(to_unsigned( 9313, 16)), --  9313 / 0x2461
    3776 => std_logic_vector(to_unsigned( 6397, 16)), --  6397 / 0x18fd
    3777 => std_logic_vector(to_unsigned( 2957, 16)), --  2957 / 0x0b8d
    3778 => std_logic_vector(to_unsigned( 7288, 16)), --  7288 / 0x1c78
    3779 => std_logic_vector(to_unsigned( 5484, 16)), --  5484 / 0x156c
    3780 => std_logic_vector(to_unsigned( 6031, 16)), --  6031 / 0x178f
    3781 => std_logic_vector(to_unsigned(10217, 16)), -- 10217 / 0x27e9 -- last item of row
    3782 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    3783 => std_logic_vector(to_unsigned(10175, 16)), -- 10175 / 0x27bf
    3784 => std_logic_vector(to_unsigned( 9009, 16)), --  9009 / 0x2331
    3785 => std_logic_vector(to_unsigned( 9889, 16)), --  9889 / 0x26a1
    3786 => std_logic_vector(to_unsigned( 3091, 16)), --  3091 / 0x0c13
    3787 => std_logic_vector(to_unsigned( 4985, 16)), --  4985 / 0x1379
    3788 => std_logic_vector(to_unsigned( 7267, 16)), --  7267 / 0x1c63
    3789 => std_logic_vector(to_unsigned( 4092, 16)), --  4092 / 0x0ffc
    3790 => std_logic_vector(to_unsigned( 8874, 16)), --  8874 / 0x22aa
    3791 => std_logic_vector(to_unsigned( 5671, 16)), --  5671 / 0x1627
    3792 => std_logic_vector(to_unsigned( 2777, 16)), --  2777 / 0x0ad9
    3793 => std_logic_vector(to_unsigned( 2189, 16)), --  2189 / 0x088d
    3794 => std_logic_vector(to_unsigned( 8716, 16)), --  8716 / 0x220c -- last item of row
    3795 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    3796 => std_logic_vector(to_unsigned( 9052, 16)), --  9052 / 0x235c
    3797 => std_logic_vector(to_unsigned( 4795, 16)), --  4795 / 0x12bb
    3798 => std_logic_vector(to_unsigned( 3924, 16)), --  3924 / 0x0f54
    3799 => std_logic_vector(to_unsigned( 3370, 16)), --  3370 / 0x0d2a
    3800 => std_logic_vector(to_unsigned(10058, 16)), -- 10058 / 0x274a
    3801 => std_logic_vector(to_unsigned( 1128, 16)), --  1128 / 0x0468
    3802 => std_logic_vector(to_unsigned( 9996, 16)), --  9996 / 0x270c
    3803 => std_logic_vector(to_unsigned(10165, 16)), -- 10165 / 0x27b5
    3804 => std_logic_vector(to_unsigned( 9360, 16)), --  9360 / 0x2490
    3805 => std_logic_vector(to_unsigned( 4297, 16)), --  4297 / 0x10c9
    3806 => std_logic_vector(to_unsigned(  434, 16)), --   434 / 0x01b2
    3807 => std_logic_vector(to_unsigned( 5138, 16)), --  5138 / 0x1412 -- last item of row
    3808 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    3809 => std_logic_vector(to_unsigned( 2379, 16)), --  2379 / 0x094b
    3810 => std_logic_vector(to_unsigned( 7834, 16)), --  7834 / 0x1e9a
    3811 => std_logic_vector(to_unsigned( 4835, 16)), --  4835 / 0x12e3
    3812 => std_logic_vector(to_unsigned( 2327, 16)), --  2327 / 0x0917
    3813 => std_logic_vector(to_unsigned( 9843, 16)), --  9843 / 0x2673
    3814 => std_logic_vector(to_unsigned(  804, 16)), --   804 / 0x0324
    3815 => std_logic_vector(to_unsigned(  329, 16)), --   329 / 0x0149
    3816 => std_logic_vector(to_unsigned( 8353, 16)), --  8353 / 0x20a1
    3817 => std_logic_vector(to_unsigned( 7167, 16)), --  7167 / 0x1bff
    3818 => std_logic_vector(to_unsigned( 3070, 16)), --  3070 / 0x0bfe
    3819 => std_logic_vector(to_unsigned( 1528, 16)), --  1528 / 0x05f8
    3820 => std_logic_vector(to_unsigned( 7311, 16)), --  7311 / 0x1c8f -- last item of row
    3821 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    3822 => std_logic_vector(to_unsigned( 3435, 16)), --  3435 / 0x0d6b
    3823 => std_logic_vector(to_unsigned( 7871, 16)), --  7871 / 0x1ebf
    3824 => std_logic_vector(to_unsigned(  348, 16)), --   348 / 0x015c
    3825 => std_logic_vector(to_unsigned( 3693, 16)), --  3693 / 0x0e6d
    3826 => std_logic_vector(to_unsigned( 1876, 16)), --  1876 / 0x0754
    3827 => std_logic_vector(to_unsigned( 6585, 16)), --  6585 / 0x19b9
    3828 => std_logic_vector(to_unsigned(10340, 16)), -- 10340 / 0x2864
    3829 => std_logic_vector(to_unsigned( 7144, 16)), --  7144 / 0x1be8
    3830 => std_logic_vector(to_unsigned( 5870, 16)), --  5870 / 0x16ee
    3831 => std_logic_vector(to_unsigned( 2084, 16)), --  2084 / 0x0824
    3832 => std_logic_vector(to_unsigned( 4052, 16)), --  4052 / 0x0fd4
    3833 => std_logic_vector(to_unsigned( 2780, 16)), --  2780 / 0x0adc -- last item of row
    3834 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    3835 => std_logic_vector(to_unsigned( 3917, 16)), --  3917 / 0x0f4d
    3836 => std_logic_vector(to_unsigned( 3111, 16)), --  3111 / 0x0c27
    3837 => std_logic_vector(to_unsigned( 3476, 16)), --  3476 / 0x0d94
    3838 => std_logic_vector(to_unsigned( 1304, 16)), --  1304 / 0x0518
    3839 => std_logic_vector(to_unsigned(10331, 16)), -- 10331 / 0x285b
    3840 => std_logic_vector(to_unsigned( 5939, 16)), --  5939 / 0x1733
    3841 => std_logic_vector(to_unsigned( 5199, 16)), --  5199 / 0x144f
    3842 => std_logic_vector(to_unsigned( 1611, 16)), --  1611 / 0x064b
    3843 => std_logic_vector(to_unsigned( 1991, 16)), --  1991 / 0x07c7
    3844 => std_logic_vector(to_unsigned(  699, 16)), --   699 / 0x02bb
    3845 => std_logic_vector(to_unsigned( 8316, 16)), --  8316 / 0x207c
    3846 => std_logic_vector(to_unsigned( 9960, 16)), --  9960 / 0x26e8 -- last item of row
    3847 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    3848 => std_logic_vector(to_unsigned( 6883, 16)), --  6883 / 0x1ae3
    3849 => std_logic_vector(to_unsigned( 3237, 16)), --  3237 / 0x0ca5
    3850 => std_logic_vector(to_unsigned( 1717, 16)), --  1717 / 0x06b5
    3851 => std_logic_vector(to_unsigned(10752, 16)), -- 10752 / 0x2a00
    3852 => std_logic_vector(to_unsigned( 7891, 16)), --  7891 / 0x1ed3
    3853 => std_logic_vector(to_unsigned( 9764, 16)), --  9764 / 0x2624
    3854 => std_logic_vector(to_unsigned( 4745, 16)), --  4745 / 0x1289
    3855 => std_logic_vector(to_unsigned( 3888, 16)), --  3888 / 0x0f30
    3856 => std_logic_vector(to_unsigned(10009, 16)), -- 10009 / 0x2719
    3857 => std_logic_vector(to_unsigned( 4176, 16)), --  4176 / 0x1050
    3858 => std_logic_vector(to_unsigned( 4614, 16)), --  4614 / 0x1206
    3859 => std_logic_vector(to_unsigned( 1567, 16)), --  1567 / 0x061f -- last item of row
    3860 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    3861 => std_logic_vector(to_unsigned(10587, 16)), -- 10587 / 0x295b
    3862 => std_logic_vector(to_unsigned( 2195, 16)), --  2195 / 0x0893
    3863 => std_logic_vector(to_unsigned( 1689, 16)), --  1689 / 0x0699
    3864 => std_logic_vector(to_unsigned( 2968, 16)), --  2968 / 0x0b98
    3865 => std_logic_vector(to_unsigned( 5420, 16)), --  5420 / 0x152c
    3866 => std_logic_vector(to_unsigned( 2580, 16)), --  2580 / 0x0a14
    3867 => std_logic_vector(to_unsigned( 2883, 16)), --  2883 / 0x0b43
    3868 => std_logic_vector(to_unsigned( 6496, 16)), --  6496 / 0x1960
    3869 => std_logic_vector(to_unsigned(  111, 16)), --   111 / 0x006f
    3870 => std_logic_vector(to_unsigned( 6023, 16)), --  6023 / 0x1787
    3871 => std_logic_vector(to_unsigned( 1024, 16)), --  1024 / 0x0400
    3872 => std_logic_vector(to_unsigned( 4449, 16)), --  4449 / 0x1161 -- last item of row
    3873 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    3874 => std_logic_vector(to_unsigned( 3786, 16)), --  3786 / 0x0eca
    3875 => std_logic_vector(to_unsigned( 8593, 16)), --  8593 / 0x2191
    3876 => std_logic_vector(to_unsigned( 2074, 16)), --  2074 / 0x081a
    3877 => std_logic_vector(to_unsigned( 3321, 16)), --  3321 / 0x0cf9
    3878 => std_logic_vector(to_unsigned( 5057, 16)), --  5057 / 0x13c1
    3879 => std_logic_vector(to_unsigned( 1450, 16)), --  1450 / 0x05aa
    3880 => std_logic_vector(to_unsigned( 3840, 16)), --  3840 / 0x0f00
    3881 => std_logic_vector(to_unsigned( 5444, 16)), --  5444 / 0x1544
    3882 => std_logic_vector(to_unsigned( 6572, 16)), --  6572 / 0x19ac
    3883 => std_logic_vector(to_unsigned( 3094, 16)), --  3094 / 0x0c16
    3884 => std_logic_vector(to_unsigned( 9892, 16)), --  9892 / 0x26a4
    3885 => std_logic_vector(to_unsigned( 1512, 16)), --  1512 / 0x05e8 -- last item of row
    3886 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    3887 => std_logic_vector(to_unsigned( 8548, 16)), --  8548 / 0x2164
    3888 => std_logic_vector(to_unsigned( 1848, 16)), --  1848 / 0x0738
    3889 => std_logic_vector(to_unsigned(10372, 16)), -- 10372 / 0x2884
    3890 => std_logic_vector(to_unsigned( 4585, 16)), --  4585 / 0x11e9
    3891 => std_logic_vector(to_unsigned( 7313, 16)), --  7313 / 0x1c91
    3892 => std_logic_vector(to_unsigned( 6536, 16)), --  6536 / 0x1988
    3893 => std_logic_vector(to_unsigned( 6379, 16)), --  6379 / 0x18eb
    3894 => std_logic_vector(to_unsigned( 1766, 16)), --  1766 / 0x06e6
    3895 => std_logic_vector(to_unsigned( 9462, 16)), --  9462 / 0x24f6
    3896 => std_logic_vector(to_unsigned( 2456, 16)), --  2456 / 0x0998
    3897 => std_logic_vector(to_unsigned( 5606, 16)), --  5606 / 0x15e6
    3898 => std_logic_vector(to_unsigned( 9975, 16)), --  9975 / 0x26f7 -- last item of row
    3899 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    3900 => std_logic_vector(to_unsigned( 8204, 16)), --  8204 / 0x200c
    3901 => std_logic_vector(to_unsigned(10593, 16)), -- 10593 / 0x2961
    3902 => std_logic_vector(to_unsigned( 7935, 16)), --  7935 / 0x1eff
    3903 => std_logic_vector(to_unsigned( 3636, 16)), --  3636 / 0x0e34
    3904 => std_logic_vector(to_unsigned( 3882, 16)), --  3882 / 0x0f2a
    3905 => std_logic_vector(to_unsigned(  394, 16)), --   394 / 0x018a
    3906 => std_logic_vector(to_unsigned( 5968, 16)), --  5968 / 0x1750
    3907 => std_logic_vector(to_unsigned( 8561, 16)), --  8561 / 0x2171
    3908 => std_logic_vector(to_unsigned( 2395, 16)), --  2395 / 0x095b
    3909 => std_logic_vector(to_unsigned( 7289, 16)), --  7289 / 0x1c79
    3910 => std_logic_vector(to_unsigned( 9267, 16)), --  9267 / 0x2433
    3911 => std_logic_vector(to_unsigned( 9978, 16)), --  9978 / 0x26fa -- last item of row
    3912 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    3913 => std_logic_vector(to_unsigned( 7795, 16)), --  7795 / 0x1e73
    3914 => std_logic_vector(to_unsigned(   74, 16)), --    74 / 0x004a
    3915 => std_logic_vector(to_unsigned( 1633, 16)), --  1633 / 0x0661
    3916 => std_logic_vector(to_unsigned( 9542, 16)), --  9542 / 0x2546
    3917 => std_logic_vector(to_unsigned( 6867, 16)), --  6867 / 0x1ad3
    3918 => std_logic_vector(to_unsigned( 7352, 16)), --  7352 / 0x1cb8
    3919 => std_logic_vector(to_unsigned( 6417, 16)), --  6417 / 0x1911
    3920 => std_logic_vector(to_unsigned( 7568, 16)), --  7568 / 0x1d90
    3921 => std_logic_vector(to_unsigned(10623, 16)), -- 10623 / 0x297f
    3922 => std_logic_vector(to_unsigned(  725, 16)), --   725 / 0x02d5
    3923 => std_logic_vector(to_unsigned( 2531, 16)), --  2531 / 0x09e3
    3924 => std_logic_vector(to_unsigned( 9115, 16)), --  9115 / 0x239b -- last item of row
    3925 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    3926 => std_logic_vector(to_unsigned( 7151, 16)), --  7151 / 0x1bef
    3927 => std_logic_vector(to_unsigned( 2482, 16)), --  2482 / 0x09b2
    3928 => std_logic_vector(to_unsigned( 4260, 16)), --  4260 / 0x10a4
    3929 => std_logic_vector(to_unsigned( 5003, 16)), --  5003 / 0x138b
    3930 => std_logic_vector(to_unsigned(10105, 16)), -- 10105 / 0x2779
    3931 => std_logic_vector(to_unsigned( 7419, 16)), --  7419 / 0x1cfb
    3932 => std_logic_vector(to_unsigned( 9203, 16)), --  9203 / 0x23f3
    3933 => std_logic_vector(to_unsigned( 6691, 16)), --  6691 / 0x1a23
    3934 => std_logic_vector(to_unsigned( 8798, 16)), --  8798 / 0x225e
    3935 => std_logic_vector(to_unsigned( 2092, 16)), --  2092 / 0x082c
    3936 => std_logic_vector(to_unsigned( 8263, 16)), --  8263 / 0x2047
    3937 => std_logic_vector(to_unsigned( 3755, 16)), --  3755 / 0x0eab -- last item of row
    3938 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    3939 => std_logic_vector(to_unsigned( 3600, 16)), --  3600 / 0x0e10
    3940 => std_logic_vector(to_unsigned(  570, 16)), --   570 / 0x023a
    3941 => std_logic_vector(to_unsigned( 4527, 16)), --  4527 / 0x11af
    3942 => std_logic_vector(to_unsigned(  200, 16)), --   200 / 0x00c8
    3943 => std_logic_vector(to_unsigned( 9718, 16)), --  9718 / 0x25f6
    3944 => std_logic_vector(to_unsigned( 6771, 16)), --  6771 / 0x1a73
    3945 => std_logic_vector(to_unsigned( 1995, 16)), --  1995 / 0x07cb
    3946 => std_logic_vector(to_unsigned( 8902, 16)), --  8902 / 0x22c6
    3947 => std_logic_vector(to_unsigned( 5446, 16)), --  5446 / 0x1546
    3948 => std_logic_vector(to_unsigned(  768, 16)), --   768 / 0x0300
    3949 => std_logic_vector(to_unsigned( 1103, 16)), --  1103 / 0x044f
    3950 => std_logic_vector(to_unsigned( 6520, 16)), --  6520 / 0x1978 -- last item of row
    3951 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    3952 => std_logic_vector(to_unsigned( 6304, 16)), --  6304 / 0x18a0
    3953 => std_logic_vector(to_unsigned( 7621, 16)), --  7621 / 0x1dc5 -- last item of row
    3954 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    3955 => std_logic_vector(to_unsigned( 6498, 16)), --  6498 / 0x1962
    3956 => std_logic_vector(to_unsigned( 9209, 16)), --  9209 / 0x23f9 -- last item of row
    3957 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    3958 => std_logic_vector(to_unsigned( 7293, 16)), --  7293 / 0x1c7d
    3959 => std_logic_vector(to_unsigned( 6786, 16)), --  6786 / 0x1a82 -- last item of row
    3960 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    3961 => std_logic_vector(to_unsigned( 5950, 16)), --  5950 / 0x173e
    3962 => std_logic_vector(to_unsigned( 1708, 16)), --  1708 / 0x06ac -- last item of row
    3963 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    3964 => std_logic_vector(to_unsigned( 8521, 16)), --  8521 / 0x2149
    3965 => std_logic_vector(to_unsigned( 1793, 16)), --  1793 / 0x0701 -- last item of row
    3966 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    3967 => std_logic_vector(to_unsigned( 6174, 16)), --  6174 / 0x181e
    3968 => std_logic_vector(to_unsigned( 7854, 16)), --  7854 / 0x1eae -- last item of row
    3969 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    3970 => std_logic_vector(to_unsigned( 9773, 16)), --  9773 / 0x262d
    3971 => std_logic_vector(to_unsigned( 1190, 16)), --  1190 / 0x04a6 -- last item of row
    3972 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    3973 => std_logic_vector(to_unsigned( 9517, 16)), --  9517 / 0x252d
    3974 => std_logic_vector(to_unsigned(10268, 16)), -- 10268 / 0x281c -- last item of row
    3975 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    3976 => std_logic_vector(to_unsigned( 2181, 16)), --  2181 / 0x0885
    3977 => std_logic_vector(to_unsigned( 9349, 16)), --  9349 / 0x2485 -- last item of row
    3978 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    3979 => std_logic_vector(to_unsigned( 1949, 16)), --  1949 / 0x079d
    3980 => std_logic_vector(to_unsigned( 5560, 16)), --  5560 / 0x15b8 -- last item of row
    3981 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    3982 => std_logic_vector(to_unsigned( 1556, 16)), --  1556 / 0x0614
    3983 => std_logic_vector(to_unsigned(  555, 16)), --   555 / 0x022b -- last item of row
    3984 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    3985 => std_logic_vector(to_unsigned( 8600, 16)), --  8600 / 0x2198
    3986 => std_logic_vector(to_unsigned( 3827, 16)), --  3827 / 0x0ef3 -- last item of row
    3987 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    3988 => std_logic_vector(to_unsigned( 5072, 16)), --  5072 / 0x13d0
    3989 => std_logic_vector(to_unsigned( 1057, 16)), --  1057 / 0x0421 -- last item of row
    3990 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    3991 => std_logic_vector(to_unsigned( 7928, 16)), --  7928 / 0x1ef8
    3992 => std_logic_vector(to_unsigned( 3542, 16)), --  3542 / 0x0dd6 -- last item of row
    3993 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    3994 => std_logic_vector(to_unsigned( 3226, 16)), --  3226 / 0x0c9a
    3995 => std_logic_vector(to_unsigned( 3762, 16)), --  3762 / 0x0eb2 -- last item of row
    3996 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    3997 => std_logic_vector(to_unsigned( 7045, 16)), --  7045 / 0x1b85
    3998 => std_logic_vector(to_unsigned( 2420, 16)), --  2420 / 0x0974 -- last item of row
    3999 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4000 => std_logic_vector(to_unsigned( 9645, 16)), --  9645 / 0x25ad
    4001 => std_logic_vector(to_unsigned( 2641, 16)), --  2641 / 0x0a51 -- last item of row
    4002 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4003 => std_logic_vector(to_unsigned( 2774, 16)), --  2774 / 0x0ad6
    4004 => std_logic_vector(to_unsigned( 2452, 16)), --  2452 / 0x0994 -- last item of row
    4005 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4006 => std_logic_vector(to_unsigned( 5331, 16)), --  5331 / 0x14d3
    4007 => std_logic_vector(to_unsigned( 2031, 16)), --  2031 / 0x07ef -- last item of row
    4008 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4009 => std_logic_vector(to_unsigned( 9400, 16)), --  9400 / 0x24b8
    4010 => std_logic_vector(to_unsigned( 7503, 16)), --  7503 / 0x1d4f -- last item of row
    4011 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4012 => std_logic_vector(to_unsigned( 1850, 16)), --  1850 / 0x073a
    4013 => std_logic_vector(to_unsigned( 2338, 16)), --  2338 / 0x0922 -- last item of row
    4014 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4015 => std_logic_vector(to_unsigned(10456, 16)), -- 10456 / 0x28d8
    4016 => std_logic_vector(to_unsigned( 9774, 16)), --  9774 / 0x262e -- last item of row
    4017 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4018 => std_logic_vector(to_unsigned( 1692, 16)), --  1692 / 0x069c
    4019 => std_logic_vector(to_unsigned( 9276, 16)), --  9276 / 0x243c -- last item of row
    4020 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4021 => std_logic_vector(to_unsigned(10037, 16)), -- 10037 / 0x2735
    4022 => std_logic_vector(to_unsigned( 4038, 16)), --  4038 / 0x0fc6 -- last item of row
    4023 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4024 => std_logic_vector(to_unsigned( 3964, 16)), --  3964 / 0x0f7c
    4025 => std_logic_vector(to_unsigned(  338, 16)), --   338 / 0x0152 -- last item of row
    4026 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4027 => std_logic_vector(to_unsigned( 2640, 16)), --  2640 / 0x0a50
    4028 => std_logic_vector(to_unsigned( 5087, 16)), --  5087 / 0x13df -- last item of row
    4029 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4030 => std_logic_vector(to_unsigned(  858, 16)), --   858 / 0x035a
    4031 => std_logic_vector(to_unsigned( 3473, 16)), --  3473 / 0x0d91 -- last item of row
    4032 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4033 => std_logic_vector(to_unsigned( 5582, 16)), --  5582 / 0x15ce
    4034 => std_logic_vector(to_unsigned( 5683, 16)), --  5683 / 0x1633 -- last item of row
    4035 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4036 => std_logic_vector(to_unsigned( 9523, 16)), --  9523 / 0x2533
    4037 => std_logic_vector(to_unsigned(  916, 16)), --   916 / 0x0394 -- last item of row
    4038 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4039 => std_logic_vector(to_unsigned( 4107, 16)), --  4107 / 0x100b
    4040 => std_logic_vector(to_unsigned( 1559, 16)), --  1559 / 0x0617 -- last item of row
    4041 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4042 => std_logic_vector(to_unsigned( 4506, 16)), --  4506 / 0x119a
    4043 => std_logic_vector(to_unsigned( 3491, 16)), --  3491 / 0x0da3 -- last item of row
    4044 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4045 => std_logic_vector(to_unsigned( 8191, 16)), --  8191 / 0x1fff
    4046 => std_logic_vector(to_unsigned( 4182, 16)), --  4182 / 0x1056 -- last item of row
    4047 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4048 => std_logic_vector(to_unsigned(10192, 16)), -- 10192 / 0x27d0
    4049 => std_logic_vector(to_unsigned( 6157, 16)), --  6157 / 0x180d -- last item of row
    4050 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4051 => std_logic_vector(to_unsigned( 5668, 16)), --  5668 / 0x1624
    4052 => std_logic_vector(to_unsigned( 3305, 16)), --  3305 / 0x0ce9 -- last item of row
    4053 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4054 => std_logic_vector(to_unsigned( 3449, 16)), --  3449 / 0x0d79
    4055 => std_logic_vector(to_unsigned( 1540, 16)), --  1540 / 0x0604 -- last item of row
    4056 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    4057 => std_logic_vector(to_unsigned( 4766, 16)), --  4766 / 0x129e
    4058 => std_logic_vector(to_unsigned( 2697, 16)), --  2697 / 0x0a89 -- last item of row
    4059 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    4060 => std_logic_vector(to_unsigned( 4069, 16)), --  4069 / 0x0fe5
    4061 => std_logic_vector(to_unsigned( 6675, 16)), --  6675 / 0x1a13 -- last item of row
    4062 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    4063 => std_logic_vector(to_unsigned( 1117, 16)), --  1117 / 0x045d
    4064 => std_logic_vector(to_unsigned( 1016, 16)), --  1016 / 0x03f8 -- last item of row
    4065 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    4066 => std_logic_vector(to_unsigned( 5619, 16)), --  5619 / 0x15f3
    4067 => std_logic_vector(to_unsigned( 3085, 16)), --  3085 / 0x0c0d -- last item of row
    4068 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    4069 => std_logic_vector(to_unsigned( 8483, 16)), --  8483 / 0x2123
    4070 => std_logic_vector(to_unsigned( 8400, 16)), --  8400 / 0x20d0 -- last item of row
    4071 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    4072 => std_logic_vector(to_unsigned( 8255, 16)), --  8255 / 0x203f
    4073 => std_logic_vector(to_unsigned(  394, 16)), --   394 / 0x018a -- last item of row
    4074 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    4075 => std_logic_vector(to_unsigned( 6338, 16)), --  6338 / 0x18c2
    4076 => std_logic_vector(to_unsigned( 5042, 16)), --  5042 / 0x13b2 -- last item of row
    4077 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    4078 => std_logic_vector(to_unsigned( 6174, 16)), --  6174 / 0x181e
    4079 => std_logic_vector(to_unsigned( 5119, 16)), --  5119 / 0x13ff -- last item of row
    4080 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    4081 => std_logic_vector(to_unsigned( 7203, 16)), --  7203 / 0x1c23
    4082 => std_logic_vector(to_unsigned( 1989, 16)), --  1989 / 0x07c5 -- last item of row
    4083 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    4084 => std_logic_vector(to_unsigned( 1781, 16)), --  1781 / 0x06f5
    4085 => std_logic_vector(to_unsigned( 5174, 16)), --  5174 / 0x1436 -- last item of row
    4086 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4087 => std_logic_vector(to_unsigned( 1464, 16)), --  1464 / 0x05b8
    4088 => std_logic_vector(to_unsigned( 3559, 16)), --  3559 / 0x0de7 -- last item of row
    4089 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4090 => std_logic_vector(to_unsigned( 3376, 16)), --  3376 / 0x0d30
    4091 => std_logic_vector(to_unsigned( 4214, 16)), --  4214 / 0x1076 -- last item of row
    4092 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4093 => std_logic_vector(to_unsigned( 7238, 16)), --  7238 / 0x1c46
    4094 => std_logic_vector(to_unsigned(   67, 16)), --    67 / 0x0043 -- last item of row
    4095 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4096 => std_logic_vector(to_unsigned(10595, 16)), -- 10595 / 0x2963
    4097 => std_logic_vector(to_unsigned( 8831, 16)), --  8831 / 0x227f -- last item of row
    4098 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4099 => std_logic_vector(to_unsigned( 1221, 16)), --  1221 / 0x04c5
    4100 => std_logic_vector(to_unsigned( 6513, 16)), --  6513 / 0x1971 -- last item of row
    4101 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4102 => std_logic_vector(to_unsigned( 5300, 16)), --  5300 / 0x14b4
    4103 => std_logic_vector(to_unsigned( 4652, 16)), --  4652 / 0x122c -- last item of row
    4104 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4105 => std_logic_vector(to_unsigned( 1429, 16)), --  1429 / 0x0595
    4106 => std_logic_vector(to_unsigned( 9749, 16)), --  9749 / 0x2615 -- last item of row
    4107 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4108 => std_logic_vector(to_unsigned( 7878, 16)), --  7878 / 0x1ec6
    4109 => std_logic_vector(to_unsigned( 5131, 16)), --  5131 / 0x140b -- last item of row
    4110 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4111 => std_logic_vector(to_unsigned( 4435, 16)), --  4435 / 0x1153
    4112 => std_logic_vector(to_unsigned(10284, 16)), -- 10284 / 0x282c -- last item of row
    4113 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4114 => std_logic_vector(to_unsigned( 6331, 16)), --  6331 / 0x18bb
    4115 => std_logic_vector(to_unsigned( 5507, 16)), --  5507 / 0x1583 -- last item of row
    4116 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4117 => std_logic_vector(to_unsigned( 6662, 16)), --  6662 / 0x1a06
    4118 => std_logic_vector(to_unsigned( 4941, 16)), --  4941 / 0x134d -- last item of row
    4119 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4120 => std_logic_vector(to_unsigned( 9614, 16)), --  9614 / 0x258e
    4121 => std_logic_vector(to_unsigned(10238, 16)), -- 10238 / 0x27fe -- last item of row
    4122 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4123 => std_logic_vector(to_unsigned( 8400, 16)), --  8400 / 0x20d0
    4124 => std_logic_vector(to_unsigned( 8025, 16)), --  8025 / 0x1f59 -- last item of row
    4125 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4126 => std_logic_vector(to_unsigned( 9156, 16)), --  9156 / 0x23c4
    4127 => std_logic_vector(to_unsigned( 5630, 16)), --  5630 / 0x15fe -- last item of row
    4128 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4129 => std_logic_vector(to_unsigned( 7067, 16)), --  7067 / 0x1b9b
    4130 => std_logic_vector(to_unsigned( 8878, 16)), --  8878 / 0x22ae -- last item of row
    4131 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4132 => std_logic_vector(to_unsigned( 9027, 16)), --  9027 / 0x2343
    4133 => std_logic_vector(to_unsigned( 3415, 16)), --  3415 / 0x0d57 -- last item of row
    4134 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4135 => std_logic_vector(to_unsigned( 1690, 16)), --  1690 / 0x069a
    4136 => std_logic_vector(to_unsigned( 3866, 16)), --  3866 / 0x0f1a -- last item of row
    4137 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4138 => std_logic_vector(to_unsigned( 2854, 16)), --  2854 / 0x0b26
    4139 => std_logic_vector(to_unsigned( 8469, 16)), --  8469 / 0x2115 -- last item of row
    4140 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4141 => std_logic_vector(to_unsigned( 6206, 16)), --  6206 / 0x183e
    4142 => std_logic_vector(to_unsigned(  630, 16)), --   630 / 0x0276 -- last item of row
    4143 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4144 => std_logic_vector(to_unsigned(  363, 16)), --   363 / 0x016b
    4145 => std_logic_vector(to_unsigned( 5453, 16)), --  5453 / 0x154d -- last item of row
    4146 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    4147 => std_logic_vector(to_unsigned( 4125, 16)), --  4125 / 0x101d
    4148 => std_logic_vector(to_unsigned( 7008, 16)), --  7008 / 0x1b60 -- last item of row
    4149 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    4150 => std_logic_vector(to_unsigned( 1612, 16)), --  1612 / 0x064c
    4151 => std_logic_vector(to_unsigned( 6702, 16)), --  6702 / 0x1a2e -- last item of row
    4152 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    4153 => std_logic_vector(to_unsigned( 9069, 16)), --  9069 / 0x236d
    4154 => std_logic_vector(to_unsigned( 9226, 16)), --  9226 / 0x240a -- last item of row
    4155 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    4156 => std_logic_vector(to_unsigned( 5767, 16)), --  5767 / 0x1687
    4157 => std_logic_vector(to_unsigned( 4060, 16)), --  4060 / 0x0fdc -- last item of row
    4158 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    4159 => std_logic_vector(to_unsigned( 3743, 16)), --  3743 / 0x0e9f
    4160 => std_logic_vector(to_unsigned( 9237, 16)), --  9237 / 0x2415 -- last item of row
    4161 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    4162 => std_logic_vector(to_unsigned( 7018, 16)), --  7018 / 0x1b6a
    4163 => std_logic_vector(to_unsigned( 5572, 16)), --  5572 / 0x15c4 -- last item of row
    4164 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    4165 => std_logic_vector(to_unsigned( 8892, 16)), --  8892 / 0x22bc
    4166 => std_logic_vector(to_unsigned( 4536, 16)), --  4536 / 0x11b8 -- last item of row
    4167 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    4168 => std_logic_vector(to_unsigned(  853, 16)), --   853 / 0x0355
    4169 => std_logic_vector(to_unsigned( 6064, 16)), --  6064 / 0x17b0 -- last item of row
    4170 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    4171 => std_logic_vector(to_unsigned( 8069, 16)), --  8069 / 0x1f85
    4172 => std_logic_vector(to_unsigned( 5893, 16)), --  5893 / 0x1705 -- last item of row
    4173 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    4174 => std_logic_vector(to_unsigned( 2051, 16)), --  2051 / 0x0803
    4175 => std_logic_vector(to_unsigned( 2885, 16)), --  2885 / 0x0b45 -- last item of row
    4176 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4177 => std_logic_vector(to_unsigned(10691, 16)), -- 10691 / 0x29c3
    4178 => std_logic_vector(to_unsigned( 3153, 16)), --  3153 / 0x0c51 -- last item of row
    4179 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4180 => std_logic_vector(to_unsigned( 3602, 16)), --  3602 / 0x0e12
    4181 => std_logic_vector(to_unsigned( 4055, 16)), --  4055 / 0x0fd7 -- last item of row
    4182 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4183 => std_logic_vector(to_unsigned(  328, 16)), --   328 / 0x0148
    4184 => std_logic_vector(to_unsigned( 1717, 16)), --  1717 / 0x06b5 -- last item of row
    4185 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4186 => std_logic_vector(to_unsigned( 2219, 16)), --  2219 / 0x08ab
    4187 => std_logic_vector(to_unsigned( 9299, 16)), --  9299 / 0x2453 -- last item of row
    4188 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4189 => std_logic_vector(to_unsigned( 1939, 16)), --  1939 / 0x0793
    4190 => std_logic_vector(to_unsigned( 7898, 16)), --  7898 / 0x1eda -- last item of row
    4191 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4192 => std_logic_vector(to_unsigned(  617, 16)), --   617 / 0x0269
    4193 => std_logic_vector(to_unsigned(  206, 16)), --   206 / 0x00ce -- last item of row
    4194 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4195 => std_logic_vector(to_unsigned( 8544, 16)), --  8544 / 0x2160
    4196 => std_logic_vector(to_unsigned( 1374, 16)), --  1374 / 0x055e -- last item of row
    4197 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4198 => std_logic_vector(to_unsigned(10676, 16)), -- 10676 / 0x29b4
    4199 => std_logic_vector(to_unsigned( 3240, 16)), --  3240 / 0x0ca8 -- last item of row
    4200 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4201 => std_logic_vector(to_unsigned( 6672, 16)), --  6672 / 0x1a10
    4202 => std_logic_vector(to_unsigned( 9489, 16)), --  9489 / 0x2511 -- last item of row
    4203 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4204 => std_logic_vector(to_unsigned( 3170, 16)), --  3170 / 0x0c62
    4205 => std_logic_vector(to_unsigned( 7457, 16)), --  7457 / 0x1d21 -- last item of row
    4206 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4207 => std_logic_vector(to_unsigned( 7868, 16)), --  7868 / 0x1ebc
    4208 => std_logic_vector(to_unsigned( 5731, 16)), --  5731 / 0x1663 -- last item of row
    4209 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4210 => std_logic_vector(to_unsigned( 6121, 16)), --  6121 / 0x17e9
    4211 => std_logic_vector(to_unsigned(10732, 16)), -- 10732 / 0x29ec -- last item of row
    4212 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4213 => std_logic_vector(to_unsigned( 4843, 16)), --  4843 / 0x12eb
    4214 => std_logic_vector(to_unsigned( 9132, 16)), --  9132 / 0x23ac -- last item of row
    4215 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4216 => std_logic_vector(to_unsigned(  580, 16)), --   580 / 0x0244
    4217 => std_logic_vector(to_unsigned( 9591, 16)), --  9591 / 0x2577 -- last item of row
    4218 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4219 => std_logic_vector(to_unsigned( 6267, 16)), --  6267 / 0x187b
    4220 => std_logic_vector(to_unsigned( 9290, 16)), --  9290 / 0x244a -- last item of row
    4221 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4222 => std_logic_vector(to_unsigned( 3009, 16)), --  3009 / 0x0bc1
    4223 => std_logic_vector(to_unsigned( 2268, 16)), --  2268 / 0x08dc -- last item of row
    4224 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4225 => std_logic_vector(to_unsigned(  195, 16)), --   195 / 0x00c3
    4226 => std_logic_vector(to_unsigned( 2419, 16)), --  2419 / 0x0973 -- last item of row
    4227 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4228 => std_logic_vector(to_unsigned( 8016, 16)), --  8016 / 0x1f50
    4229 => std_logic_vector(to_unsigned( 1557, 16)), --  1557 / 0x0615 -- last item of row
    4230 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4231 => std_logic_vector(to_unsigned( 1516, 16)), --  1516 / 0x05ec
    4232 => std_logic_vector(to_unsigned( 9195, 16)), --  9195 / 0x23eb -- last item of row
    4233 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4234 => std_logic_vector(to_unsigned( 8062, 16)), --  8062 / 0x1f7e
    4235 => std_logic_vector(to_unsigned( 9064, 16)), --  9064 / 0x2368 -- last item of row
    4236 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    4237 => std_logic_vector(to_unsigned( 2095, 16)), --  2095 / 0x082f
    4238 => std_logic_vector(to_unsigned( 8968, 16)), --  8968 / 0x2308 -- last item of row
    4239 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    4240 => std_logic_vector(to_unsigned(  753, 16)), --   753 / 0x02f1
    4241 => std_logic_vector(to_unsigned( 7326, 16)), --  7326 / 0x1c9e -- last item of row
    4242 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    4243 => std_logic_vector(to_unsigned( 6291, 16)), --  6291 / 0x1893
    4244 => std_logic_vector(to_unsigned( 3833, 16)), --  3833 / 0x0ef9 -- last item of row
    4245 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    4246 => std_logic_vector(to_unsigned( 2614, 16)), --  2614 / 0x0a36
    4247 => std_logic_vector(to_unsigned( 7844, 16)), --  7844 / 0x1ea4 -- last item of row
    4248 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    4249 => std_logic_vector(to_unsigned( 2303, 16)), --  2303 / 0x08ff
    4250 => std_logic_vector(to_unsigned(  646, 16)), --   646 / 0x0286 -- last item of row
    4251 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    4252 => std_logic_vector(to_unsigned( 2075, 16)), --  2075 / 0x081b
    4253 => std_logic_vector(to_unsigned(  611, 16)), --   611 / 0x0263 -- last item of row
    4254 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    4255 => std_logic_vector(to_unsigned( 4687, 16)), --  4687 / 0x124f
    4256 => std_logic_vector(to_unsigned(  362, 16)), --   362 / 0x016a -- last item of row
    4257 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    4258 => std_logic_vector(to_unsigned( 8684, 16)), --  8684 / 0x21ec
    4259 => std_logic_vector(to_unsigned( 9940, 16)), --  9940 / 0x26d4 -- last item of row
    4260 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    4261 => std_logic_vector(to_unsigned( 4830, 16)), --  4830 / 0x12de
    4262 => std_logic_vector(to_unsigned( 2065, 16)), --  2065 / 0x0811 -- last item of row
    4263 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    4264 => std_logic_vector(to_unsigned( 7038, 16)), --  7038 / 0x1b7e
    4265 => std_logic_vector(to_unsigned( 1363, 16)), --  1363 / 0x0553 -- last item of row
    4266 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4267 => std_logic_vector(to_unsigned( 1769, 16)), --  1769 / 0x06e9
    4268 => std_logic_vector(to_unsigned( 7837, 16)), --  7837 / 0x1e9d -- last item of row
    4269 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4270 => std_logic_vector(to_unsigned( 3801, 16)), --  3801 / 0x0ed9
    4271 => std_logic_vector(to_unsigned( 1689, 16)), --  1689 / 0x0699 -- last item of row
    4272 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4273 => std_logic_vector(to_unsigned(10070, 16)), -- 10070 / 0x2756
    4274 => std_logic_vector(to_unsigned( 2359, 16)), --  2359 / 0x0937 -- last item of row
    4275 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4276 => std_logic_vector(to_unsigned( 3667, 16)), --  3667 / 0x0e53
    4277 => std_logic_vector(to_unsigned( 9918, 16)), --  9918 / 0x26be -- last item of row
    4278 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4279 => std_logic_vector(to_unsigned( 1914, 16)), --  1914 / 0x077a
    4280 => std_logic_vector(to_unsigned( 6920, 16)), --  6920 / 0x1b08 -- last item of row
    4281 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4282 => std_logic_vector(to_unsigned( 4244, 16)), --  4244 / 0x1094
    4283 => std_logic_vector(to_unsigned( 5669, 16)), --  5669 / 0x1625 -- last item of row
    4284 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4285 => std_logic_vector(to_unsigned(10245, 16)), -- 10245 / 0x2805
    4286 => std_logic_vector(to_unsigned( 7821, 16)), --  7821 / 0x1e8d -- last item of row
    4287 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4288 => std_logic_vector(to_unsigned( 7648, 16)), --  7648 / 0x1de0
    4289 => std_logic_vector(to_unsigned( 3944, 16)), --  3944 / 0x0f68 -- last item of row
    4290 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4291 => std_logic_vector(to_unsigned( 3310, 16)), --  3310 / 0x0cee
    4292 => std_logic_vector(to_unsigned( 5488, 16)), --  5488 / 0x1570 -- last item of row
    4293 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4294 => std_logic_vector(to_unsigned( 6346, 16)), --  6346 / 0x18ca
    4295 => std_logic_vector(to_unsigned( 9666, 16)), --  9666 / 0x25c2 -- last item of row
    4296 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4297 => std_logic_vector(to_unsigned( 7088, 16)), --  7088 / 0x1bb0
    4298 => std_logic_vector(to_unsigned( 6122, 16)), --  6122 / 0x17ea -- last item of row
    4299 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4300 => std_logic_vector(to_unsigned( 1291, 16)), --  1291 / 0x050b
    4301 => std_logic_vector(to_unsigned( 7827, 16)), --  7827 / 0x1e93 -- last item of row
    4302 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4303 => std_logic_vector(to_unsigned(10592, 16)), -- 10592 / 0x2960
    4304 => std_logic_vector(to_unsigned( 8945, 16)), --  8945 / 0x22f1 -- last item of row
    4305 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4306 => std_logic_vector(to_unsigned( 3609, 16)), --  3609 / 0x0e19
    4307 => std_logic_vector(to_unsigned( 7120, 16)), --  7120 / 0x1bd0 -- last item of row
    4308 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4309 => std_logic_vector(to_unsigned( 9168, 16)), --  9168 / 0x23d0
    4310 => std_logic_vector(to_unsigned( 9112, 16)), --  9112 / 0x2398 -- last item of row
    4311 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4312 => std_logic_vector(to_unsigned( 6203, 16)), --  6203 / 0x183b
    4313 => std_logic_vector(to_unsigned( 8052, 16)), --  8052 / 0x1f74 -- last item of row
    4314 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4315 => std_logic_vector(to_unsigned( 3330, 16)), --  3330 / 0x0d02
    4316 => std_logic_vector(to_unsigned( 2895, 16)), --  2895 / 0x0b4f -- last item of row
    4317 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4318 => std_logic_vector(to_unsigned( 4264, 16)), --  4264 / 0x10a8
    4319 => std_logic_vector(to_unsigned(10563, 16)), -- 10563 / 0x2943 -- last item of row
    4320 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4321 => std_logic_vector(to_unsigned(10556, 16)), -- 10556 / 0x293c
    4322 => std_logic_vector(to_unsigned( 6496, 16)), --  6496 / 0x1960 -- last item of row
    4323 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4324 => std_logic_vector(to_unsigned( 8807, 16)), --  8807 / 0x2267
    4325 => std_logic_vector(to_unsigned( 7645, 16)), --  7645 / 0x1ddd -- last item of row
    4326 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    4327 => std_logic_vector(to_unsigned( 1999, 16)), --  1999 / 0x07cf
    4328 => std_logic_vector(to_unsigned( 4530, 16)), --  4530 / 0x11b2 -- last item of row
    4329 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    4330 => std_logic_vector(to_unsigned( 9202, 16)), --  9202 / 0x23f2
    4331 => std_logic_vector(to_unsigned( 6818, 16)), --  6818 / 0x1aa2 -- last item of row
    4332 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    4333 => std_logic_vector(to_unsigned( 3403, 16)), --  3403 / 0x0d4b
    4334 => std_logic_vector(to_unsigned( 1734, 16)), --  1734 / 0x06c6 -- last item of row
    4335 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    4336 => std_logic_vector(to_unsigned( 2106, 16)), --  2106 / 0x083a
    4337 => std_logic_vector(to_unsigned( 9023, 16)), --  9023 / 0x233f -- last item of row
    4338 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    4339 => std_logic_vector(to_unsigned( 6881, 16)), --  6881 / 0x1ae1
    4340 => std_logic_vector(to_unsigned( 3883, 16)), --  3883 / 0x0f2b -- last item of row
    4341 => std_logic_vector(to_unsigned(   25, 16)), --    25 / 0x0019
    4342 => std_logic_vector(to_unsigned( 3895, 16)), --  3895 / 0x0f37
    4343 => std_logic_vector(to_unsigned( 2171, 16)), --  2171 / 0x087b -- last item of row
    4344 => std_logic_vector(to_unsigned(   26, 16)), --    26 / 0x001a
    4345 => std_logic_vector(to_unsigned( 4062, 16)), --  4062 / 0x0fde
    4346 => std_logic_vector(to_unsigned( 6424, 16)), --  6424 / 0x1918 -- last item of row
    4347 => std_logic_vector(to_unsigned(   27, 16)), --    27 / 0x001b
    4348 => std_logic_vector(to_unsigned( 3755, 16)), --  3755 / 0x0eab
    4349 => std_logic_vector(to_unsigned( 9536, 16)), --  9536 / 0x2540 -- last item of row
    4350 => std_logic_vector(to_unsigned(   28, 16)), --    28 / 0x001c
    4351 => std_logic_vector(to_unsigned( 4683, 16)), --  4683 / 0x124b
    4352 => std_logic_vector(to_unsigned( 2131, 16)), --  2131 / 0x0853 -- last item of row
    4353 => std_logic_vector(to_unsigned(   29, 16)), --    29 / 0x001d
    4354 => std_logic_vector(to_unsigned( 7347, 16)), --  7347 / 0x1cb3
    4355 => std_logic_vector(to_unsigned( 8027, 16)), --  8027 / 0x1f5b -- last item of row
    -- Table for fecframe_normal, C8_9
    4356 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4357 => std_logic_vector(to_unsigned( 6235, 16)), --  6235 / 0x185b
    4358 => std_logic_vector(to_unsigned( 2848, 16)), --  2848 / 0x0b20
    4359 => std_logic_vector(to_unsigned( 3222, 16)), --  3222 / 0x0c96 -- last item of row
    4360 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4361 => std_logic_vector(to_unsigned( 5800, 16)), --  5800 / 0x16a8
    4362 => std_logic_vector(to_unsigned( 3492, 16)), --  3492 / 0x0da4
    4363 => std_logic_vector(to_unsigned( 5348, 16)), --  5348 / 0x14e4 -- last item of row
    4364 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4365 => std_logic_vector(to_unsigned( 2757, 16)), --  2757 / 0x0ac5
    4366 => std_logic_vector(to_unsigned(  927, 16)), --   927 / 0x039f
    4367 => std_logic_vector(to_unsigned(   90, 16)), --    90 / 0x005a -- last item of row
    4368 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4369 => std_logic_vector(to_unsigned( 6961, 16)), --  6961 / 0x1b31
    4370 => std_logic_vector(to_unsigned( 4516, 16)), --  4516 / 0x11a4
    4371 => std_logic_vector(to_unsigned( 4739, 16)), --  4739 / 0x1283 -- last item of row
    4372 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4373 => std_logic_vector(to_unsigned( 1172, 16)), --  1172 / 0x0494
    4374 => std_logic_vector(to_unsigned( 3237, 16)), --  3237 / 0x0ca5
    4375 => std_logic_vector(to_unsigned( 6264, 16)), --  6264 / 0x1878 -- last item of row
    4376 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4377 => std_logic_vector(to_unsigned( 1927, 16)), --  1927 / 0x0787
    4378 => std_logic_vector(to_unsigned( 2425, 16)), --  2425 / 0x0979
    4379 => std_logic_vector(to_unsigned( 3683, 16)), --  3683 / 0x0e63 -- last item of row
    4380 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4381 => std_logic_vector(to_unsigned( 3714, 16)), --  3714 / 0x0e82
    4382 => std_logic_vector(to_unsigned( 6309, 16)), --  6309 / 0x18a5
    4383 => std_logic_vector(to_unsigned( 2495, 16)), --  2495 / 0x09bf -- last item of row
    4384 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4385 => std_logic_vector(to_unsigned( 3070, 16)), --  3070 / 0x0bfe
    4386 => std_logic_vector(to_unsigned( 6342, 16)), --  6342 / 0x18c6
    4387 => std_logic_vector(to_unsigned( 7154, 16)), --  7154 / 0x1bf2 -- last item of row
    4388 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4389 => std_logic_vector(to_unsigned( 2428, 16)), --  2428 / 0x097c
    4390 => std_logic_vector(to_unsigned(  613, 16)), --   613 / 0x0265
    4391 => std_logic_vector(to_unsigned( 3761, 16)), --  3761 / 0x0eb1 -- last item of row
    4392 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4393 => std_logic_vector(to_unsigned( 2906, 16)), --  2906 / 0x0b5a
    4394 => std_logic_vector(to_unsigned(  264, 16)), --   264 / 0x0108
    4395 => std_logic_vector(to_unsigned( 5927, 16)), --  5927 / 0x1727 -- last item of row
    4396 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4397 => std_logic_vector(to_unsigned( 1716, 16)), --  1716 / 0x06b4
    4398 => std_logic_vector(to_unsigned( 1950, 16)), --  1950 / 0x079e
    4399 => std_logic_vector(to_unsigned( 4273, 16)), --  4273 / 0x10b1 -- last item of row
    4400 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4401 => std_logic_vector(to_unsigned( 4613, 16)), --  4613 / 0x1205
    4402 => std_logic_vector(to_unsigned( 6179, 16)), --  6179 / 0x1823
    4403 => std_logic_vector(to_unsigned( 3491, 16)), --  3491 / 0x0da3 -- last item of row
    4404 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4405 => std_logic_vector(to_unsigned( 4865, 16)), --  4865 / 0x1301
    4406 => std_logic_vector(to_unsigned( 3286, 16)), --  3286 / 0x0cd6
    4407 => std_logic_vector(to_unsigned( 6005, 16)), --  6005 / 0x1775 -- last item of row
    4408 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4409 => std_logic_vector(to_unsigned( 1343, 16)), --  1343 / 0x053f
    4410 => std_logic_vector(to_unsigned( 5923, 16)), --  5923 / 0x1723
    4411 => std_logic_vector(to_unsigned( 3529, 16)), --  3529 / 0x0dc9 -- last item of row
    4412 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4413 => std_logic_vector(to_unsigned( 4589, 16)), --  4589 / 0x11ed
    4414 => std_logic_vector(to_unsigned( 4035, 16)), --  4035 / 0x0fc3
    4415 => std_logic_vector(to_unsigned( 2132, 16)), --  2132 / 0x0854 -- last item of row
    4416 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4417 => std_logic_vector(to_unsigned( 1579, 16)), --  1579 / 0x062b
    4418 => std_logic_vector(to_unsigned( 3920, 16)), --  3920 / 0x0f50
    4419 => std_logic_vector(to_unsigned( 6737, 16)), --  6737 / 0x1a51 -- last item of row
    4420 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4421 => std_logic_vector(to_unsigned( 1644, 16)), --  1644 / 0x066c
    4422 => std_logic_vector(to_unsigned( 1191, 16)), --  1191 / 0x04a7
    4423 => std_logic_vector(to_unsigned( 5998, 16)), --  5998 / 0x176e -- last item of row
    4424 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4425 => std_logic_vector(to_unsigned( 1482, 16)), --  1482 / 0x05ca
    4426 => std_logic_vector(to_unsigned( 2381, 16)), --  2381 / 0x094d
    4427 => std_logic_vector(to_unsigned( 4620, 16)), --  4620 / 0x120c -- last item of row
    4428 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4429 => std_logic_vector(to_unsigned( 6791, 16)), --  6791 / 0x1a87
    4430 => std_logic_vector(to_unsigned( 6014, 16)), --  6014 / 0x177e
    4431 => std_logic_vector(to_unsigned( 6596, 16)), --  6596 / 0x19c4 -- last item of row
    4432 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4433 => std_logic_vector(to_unsigned( 2738, 16)), --  2738 / 0x0ab2
    4434 => std_logic_vector(to_unsigned( 5918, 16)), --  5918 / 0x171e
    4435 => std_logic_vector(to_unsigned( 3786, 16)), --  3786 / 0x0eca -- last item of row
    4436 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4437 => std_logic_vector(to_unsigned( 5156, 16)), --  5156 / 0x1424
    4438 => std_logic_vector(to_unsigned( 6166, 16)), --  6166 / 0x1816 -- last item of row
    4439 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4440 => std_logic_vector(to_unsigned( 1504, 16)), --  1504 / 0x05e0
    4441 => std_logic_vector(to_unsigned( 4356, 16)), --  4356 / 0x1104 -- last item of row
    4442 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4443 => std_logic_vector(to_unsigned(  130, 16)), --   130 / 0x0082
    4444 => std_logic_vector(to_unsigned( 1904, 16)), --  1904 / 0x0770 -- last item of row
    4445 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4446 => std_logic_vector(to_unsigned( 6027, 16)), --  6027 / 0x178b
    4447 => std_logic_vector(to_unsigned( 3187, 16)), --  3187 / 0x0c73 -- last item of row
    4448 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4449 => std_logic_vector(to_unsigned( 6718, 16)), --  6718 / 0x1a3e
    4450 => std_logic_vector(to_unsigned(  759, 16)), --   759 / 0x02f7 -- last item of row
    4451 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4452 => std_logic_vector(to_unsigned( 6240, 16)), --  6240 / 0x1860
    4453 => std_logic_vector(to_unsigned( 2870, 16)), --  2870 / 0x0b36 -- last item of row
    4454 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4455 => std_logic_vector(to_unsigned( 2343, 16)), --  2343 / 0x0927
    4456 => std_logic_vector(to_unsigned( 1311, 16)), --  1311 / 0x051f -- last item of row
    4457 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4458 => std_logic_vector(to_unsigned( 1039, 16)), --  1039 / 0x040f
    4459 => std_logic_vector(to_unsigned( 5465, 16)), --  5465 / 0x1559 -- last item of row
    4460 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4461 => std_logic_vector(to_unsigned( 6617, 16)), --  6617 / 0x19d9
    4462 => std_logic_vector(to_unsigned( 2513, 16)), --  2513 / 0x09d1 -- last item of row
    4463 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4464 => std_logic_vector(to_unsigned( 1588, 16)), --  1588 / 0x0634
    4465 => std_logic_vector(to_unsigned( 5222, 16)), --  5222 / 0x1466 -- last item of row
    4466 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4467 => std_logic_vector(to_unsigned( 6561, 16)), --  6561 / 0x19a1
    4468 => std_logic_vector(to_unsigned(  535, 16)), --   535 / 0x0217 -- last item of row
    4469 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4470 => std_logic_vector(to_unsigned( 4765, 16)), --  4765 / 0x129d
    4471 => std_logic_vector(to_unsigned( 2054, 16)), --  2054 / 0x0806 -- last item of row
    4472 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4473 => std_logic_vector(to_unsigned( 5966, 16)), --  5966 / 0x174e
    4474 => std_logic_vector(to_unsigned( 6892, 16)), --  6892 / 0x1aec -- last item of row
    4475 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4476 => std_logic_vector(to_unsigned( 1969, 16)), --  1969 / 0x07b1
    4477 => std_logic_vector(to_unsigned( 3869, 16)), --  3869 / 0x0f1d -- last item of row
    4478 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4479 => std_logic_vector(to_unsigned( 3571, 16)), --  3571 / 0x0df3
    4480 => std_logic_vector(to_unsigned( 2420, 16)), --  2420 / 0x0974 -- last item of row
    4481 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4482 => std_logic_vector(to_unsigned( 4632, 16)), --  4632 / 0x1218
    4483 => std_logic_vector(to_unsigned(  981, 16)), --   981 / 0x03d5 -- last item of row
    4484 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4485 => std_logic_vector(to_unsigned( 3215, 16)), --  3215 / 0x0c8f
    4486 => std_logic_vector(to_unsigned( 4163, 16)), --  4163 / 0x1043 -- last item of row
    4487 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4488 => std_logic_vector(to_unsigned(  973, 16)), --   973 / 0x03cd
    4489 => std_logic_vector(to_unsigned( 3117, 16)), --  3117 / 0x0c2d -- last item of row
    4490 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4491 => std_logic_vector(to_unsigned( 3802, 16)), --  3802 / 0x0eda
    4492 => std_logic_vector(to_unsigned( 6198, 16)), --  6198 / 0x1836 -- last item of row
    4493 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4494 => std_logic_vector(to_unsigned( 3794, 16)), --  3794 / 0x0ed2
    4495 => std_logic_vector(to_unsigned( 3948, 16)), --  3948 / 0x0f6c -- last item of row
    4496 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4497 => std_logic_vector(to_unsigned( 3196, 16)), --  3196 / 0x0c7c
    4498 => std_logic_vector(to_unsigned( 6126, 16)), --  6126 / 0x17ee -- last item of row
    4499 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4500 => std_logic_vector(to_unsigned(  573, 16)), --   573 / 0x023d
    4501 => std_logic_vector(to_unsigned( 1909, 16)), --  1909 / 0x0775 -- last item of row
    4502 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4503 => std_logic_vector(to_unsigned(  850, 16)), --   850 / 0x0352
    4504 => std_logic_vector(to_unsigned( 4034, 16)), --  4034 / 0x0fc2 -- last item of row
    4505 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4506 => std_logic_vector(to_unsigned( 5622, 16)), --  5622 / 0x15f6
    4507 => std_logic_vector(to_unsigned( 1601, 16)), --  1601 / 0x0641 -- last item of row
    4508 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4509 => std_logic_vector(to_unsigned( 6005, 16)), --  6005 / 0x1775
    4510 => std_logic_vector(to_unsigned(  524, 16)), --   524 / 0x020c -- last item of row
    4511 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4512 => std_logic_vector(to_unsigned( 5251, 16)), --  5251 / 0x1483
    4513 => std_logic_vector(to_unsigned( 5783, 16)), --  5783 / 0x1697 -- last item of row
    4514 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4515 => std_logic_vector(to_unsigned(  172, 16)), --   172 / 0x00ac
    4516 => std_logic_vector(to_unsigned( 2032, 16)), --  2032 / 0x07f0 -- last item of row
    4517 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4518 => std_logic_vector(to_unsigned( 1875, 16)), --  1875 / 0x0753
    4519 => std_logic_vector(to_unsigned( 2475, 16)), --  2475 / 0x09ab -- last item of row
    4520 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4521 => std_logic_vector(to_unsigned(  497, 16)), --   497 / 0x01f1
    4522 => std_logic_vector(to_unsigned( 1291, 16)), --  1291 / 0x050b -- last item of row
    4523 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4524 => std_logic_vector(to_unsigned( 2566, 16)), --  2566 / 0x0a06
    4525 => std_logic_vector(to_unsigned( 3430, 16)), --  3430 / 0x0d66 -- last item of row
    4526 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4527 => std_logic_vector(to_unsigned( 1249, 16)), --  1249 / 0x04e1
    4528 => std_logic_vector(to_unsigned(  740, 16)), --   740 / 0x02e4 -- last item of row
    4529 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4530 => std_logic_vector(to_unsigned( 2944, 16)), --  2944 / 0x0b80
    4531 => std_logic_vector(to_unsigned( 1948, 16)), --  1948 / 0x079c -- last item of row
    4532 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4533 => std_logic_vector(to_unsigned( 6528, 16)), --  6528 / 0x1980
    4534 => std_logic_vector(to_unsigned( 2899, 16)), --  2899 / 0x0b53 -- last item of row
    4535 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4536 => std_logic_vector(to_unsigned( 2243, 16)), --  2243 / 0x08c3
    4537 => std_logic_vector(to_unsigned( 3616, 16)), --  3616 / 0x0e20 -- last item of row
    4538 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4539 => std_logic_vector(to_unsigned(  867, 16)), --   867 / 0x0363
    4540 => std_logic_vector(to_unsigned( 3733, 16)), --  3733 / 0x0e95 -- last item of row
    4541 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4542 => std_logic_vector(to_unsigned( 1374, 16)), --  1374 / 0x055e
    4543 => std_logic_vector(to_unsigned( 4702, 16)), --  4702 / 0x125e -- last item of row
    4544 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4545 => std_logic_vector(to_unsigned( 4698, 16)), --  4698 / 0x125a
    4546 => std_logic_vector(to_unsigned( 2285, 16)), --  2285 / 0x08ed -- last item of row
    4547 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4548 => std_logic_vector(to_unsigned( 4760, 16)), --  4760 / 0x1298
    4549 => std_logic_vector(to_unsigned( 3917, 16)), --  3917 / 0x0f4d -- last item of row
    4550 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4551 => std_logic_vector(to_unsigned( 1859, 16)), --  1859 / 0x0743
    4552 => std_logic_vector(to_unsigned( 4058, 16)), --  4058 / 0x0fda -- last item of row
    4553 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4554 => std_logic_vector(to_unsigned( 6141, 16)), --  6141 / 0x17fd
    4555 => std_logic_vector(to_unsigned( 3527, 16)), --  3527 / 0x0dc7 -- last item of row
    4556 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4557 => std_logic_vector(to_unsigned( 2148, 16)), --  2148 / 0x0864
    4558 => std_logic_vector(to_unsigned( 5066, 16)), --  5066 / 0x13ca -- last item of row
    4559 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4560 => std_logic_vector(to_unsigned( 1306, 16)), --  1306 / 0x051a
    4561 => std_logic_vector(to_unsigned(  145, 16)), --   145 / 0x0091 -- last item of row
    4562 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4563 => std_logic_vector(to_unsigned( 2319, 16)), --  2319 / 0x090f
    4564 => std_logic_vector(to_unsigned(  871, 16)), --   871 / 0x0367 -- last item of row
    4565 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4566 => std_logic_vector(to_unsigned( 3463, 16)), --  3463 / 0x0d87
    4567 => std_logic_vector(to_unsigned( 1061, 16)), --  1061 / 0x0425 -- last item of row
    4568 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4569 => std_logic_vector(to_unsigned( 5554, 16)), --  5554 / 0x15b2
    4570 => std_logic_vector(to_unsigned( 6647, 16)), --  6647 / 0x19f7 -- last item of row
    4571 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4572 => std_logic_vector(to_unsigned( 5837, 16)), --  5837 / 0x16cd
    4573 => std_logic_vector(to_unsigned(  339, 16)), --   339 / 0x0153 -- last item of row
    4574 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4575 => std_logic_vector(to_unsigned( 5821, 16)), --  5821 / 0x16bd
    4576 => std_logic_vector(to_unsigned( 4932, 16)), --  4932 / 0x1344 -- last item of row
    4577 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4578 => std_logic_vector(to_unsigned( 6356, 16)), --  6356 / 0x18d4
    4579 => std_logic_vector(to_unsigned( 4756, 16)), --  4756 / 0x1294 -- last item of row
    4580 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4581 => std_logic_vector(to_unsigned( 3930, 16)), --  3930 / 0x0f5a
    4582 => std_logic_vector(to_unsigned(  418, 16)), --   418 / 0x01a2 -- last item of row
    4583 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4584 => std_logic_vector(to_unsigned(  211, 16)), --   211 / 0x00d3
    4585 => std_logic_vector(to_unsigned( 3094, 16)), --  3094 / 0x0c16 -- last item of row
    4586 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4587 => std_logic_vector(to_unsigned( 1007, 16)), --  1007 / 0x03ef
    4588 => std_logic_vector(to_unsigned( 4928, 16)), --  4928 / 0x1340 -- last item of row
    4589 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4590 => std_logic_vector(to_unsigned( 3584, 16)), --  3584 / 0x0e00
    4591 => std_logic_vector(to_unsigned( 1235, 16)), --  1235 / 0x04d3 -- last item of row
    4592 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4593 => std_logic_vector(to_unsigned( 6982, 16)), --  6982 / 0x1b46
    4594 => std_logic_vector(to_unsigned( 2869, 16)), --  2869 / 0x0b35 -- last item of row
    4595 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4596 => std_logic_vector(to_unsigned( 1612, 16)), --  1612 / 0x064c
    4597 => std_logic_vector(to_unsigned( 1013, 16)), --  1013 / 0x03f5 -- last item of row
    4598 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4599 => std_logic_vector(to_unsigned(  953, 16)), --   953 / 0x03b9
    4600 => std_logic_vector(to_unsigned( 4964, 16)), --  4964 / 0x1364 -- last item of row
    4601 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4602 => std_logic_vector(to_unsigned( 4555, 16)), --  4555 / 0x11cb
    4603 => std_logic_vector(to_unsigned( 4410, 16)), --  4410 / 0x113a -- last item of row
    4604 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4605 => std_logic_vector(to_unsigned( 4925, 16)), --  4925 / 0x133d
    4606 => std_logic_vector(to_unsigned( 4842, 16)), --  4842 / 0x12ea -- last item of row
    4607 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4608 => std_logic_vector(to_unsigned( 5778, 16)), --  5778 / 0x1692
    4609 => std_logic_vector(to_unsigned(  600, 16)), --   600 / 0x0258 -- last item of row
    4610 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4611 => std_logic_vector(to_unsigned( 6509, 16)), --  6509 / 0x196d
    4612 => std_logic_vector(to_unsigned( 2417, 16)), --  2417 / 0x0971 -- last item of row
    4613 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4614 => std_logic_vector(to_unsigned( 1260, 16)), --  1260 / 0x04ec
    4615 => std_logic_vector(to_unsigned( 4903, 16)), --  4903 / 0x1327 -- last item of row
    4616 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4617 => std_logic_vector(to_unsigned( 3369, 16)), --  3369 / 0x0d29
    4618 => std_logic_vector(to_unsigned( 3031, 16)), --  3031 / 0x0bd7 -- last item of row
    4619 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4620 => std_logic_vector(to_unsigned( 3557, 16)), --  3557 / 0x0de5
    4621 => std_logic_vector(to_unsigned( 3224, 16)), --  3224 / 0x0c98 -- last item of row
    4622 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4623 => std_logic_vector(to_unsigned( 3028, 16)), --  3028 / 0x0bd4
    4624 => std_logic_vector(to_unsigned(  583, 16)), --   583 / 0x0247 -- last item of row
    4625 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4626 => std_logic_vector(to_unsigned( 3258, 16)), --  3258 / 0x0cba
    4627 => std_logic_vector(to_unsigned(  440, 16)), --   440 / 0x01b8 -- last item of row
    4628 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4629 => std_logic_vector(to_unsigned( 6226, 16)), --  6226 / 0x1852
    4630 => std_logic_vector(to_unsigned( 6655, 16)), --  6655 / 0x19ff -- last item of row
    4631 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4632 => std_logic_vector(to_unsigned( 4895, 16)), --  4895 / 0x131f
    4633 => std_logic_vector(to_unsigned( 1094, 16)), --  1094 / 0x0446 -- last item of row
    4634 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4635 => std_logic_vector(to_unsigned( 1481, 16)), --  1481 / 0x05c9
    4636 => std_logic_vector(to_unsigned( 6847, 16)), --  6847 / 0x1abf -- last item of row
    4637 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4638 => std_logic_vector(to_unsigned( 4433, 16)), --  4433 / 0x1151
    4639 => std_logic_vector(to_unsigned( 1932, 16)), --  1932 / 0x078c -- last item of row
    4640 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4641 => std_logic_vector(to_unsigned( 2107, 16)), --  2107 / 0x083b
    4642 => std_logic_vector(to_unsigned( 1649, 16)), --  1649 / 0x0671 -- last item of row
    4643 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4644 => std_logic_vector(to_unsigned( 2119, 16)), --  2119 / 0x0847
    4645 => std_logic_vector(to_unsigned( 2065, 16)), --  2065 / 0x0811 -- last item of row
    4646 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4647 => std_logic_vector(to_unsigned( 4003, 16)), --  4003 / 0x0fa3
    4648 => std_logic_vector(to_unsigned( 6388, 16)), --  6388 / 0x18f4 -- last item of row
    4649 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4650 => std_logic_vector(to_unsigned( 6720, 16)), --  6720 / 0x1a40
    4651 => std_logic_vector(to_unsigned( 3622, 16)), --  3622 / 0x0e26 -- last item of row
    4652 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4653 => std_logic_vector(to_unsigned( 3694, 16)), --  3694 / 0x0e6e
    4654 => std_logic_vector(to_unsigned( 4521, 16)), --  4521 / 0x11a9 -- last item of row
    4655 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4656 => std_logic_vector(to_unsigned( 1164, 16)), --  1164 / 0x048c
    4657 => std_logic_vector(to_unsigned( 7050, 16)), --  7050 / 0x1b8a -- last item of row
    4658 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4659 => std_logic_vector(to_unsigned( 1965, 16)), --  1965 / 0x07ad
    4660 => std_logic_vector(to_unsigned( 3613, 16)), --  3613 / 0x0e1d -- last item of row
    4661 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4662 => std_logic_vector(to_unsigned( 4331, 16)), --  4331 / 0x10eb
    4663 => std_logic_vector(to_unsigned(   66, 16)), --    66 / 0x0042 -- last item of row
    4664 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4665 => std_logic_vector(to_unsigned( 2970, 16)), --  2970 / 0x0b9a
    4666 => std_logic_vector(to_unsigned( 1796, 16)), --  1796 / 0x0704 -- last item of row
    4667 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4668 => std_logic_vector(to_unsigned( 4652, 16)), --  4652 / 0x122c
    4669 => std_logic_vector(to_unsigned( 3218, 16)), --  3218 / 0x0c92 -- last item of row
    4670 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4671 => std_logic_vector(to_unsigned( 1762, 16)), --  1762 / 0x06e2
    4672 => std_logic_vector(to_unsigned( 4777, 16)), --  4777 / 0x12a9 -- last item of row
    4673 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4674 => std_logic_vector(to_unsigned( 5736, 16)), --  5736 / 0x1668
    4675 => std_logic_vector(to_unsigned( 1399, 16)), --  1399 / 0x0577 -- last item of row
    4676 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4677 => std_logic_vector(to_unsigned(  970, 16)), --   970 / 0x03ca
    4678 => std_logic_vector(to_unsigned( 2572, 16)), --  2572 / 0x0a0c -- last item of row
    4679 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4680 => std_logic_vector(to_unsigned( 2062, 16)), --  2062 / 0x080e
    4681 => std_logic_vector(to_unsigned( 6599, 16)), --  6599 / 0x19c7 -- last item of row
    4682 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4683 => std_logic_vector(to_unsigned( 4597, 16)), --  4597 / 0x11f5
    4684 => std_logic_vector(to_unsigned( 4870, 16)), --  4870 / 0x1306 -- last item of row
    4685 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4686 => std_logic_vector(to_unsigned( 1228, 16)), --  1228 / 0x04cc
    4687 => std_logic_vector(to_unsigned( 6913, 16)), --  6913 / 0x1b01 -- last item of row
    4688 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4689 => std_logic_vector(to_unsigned( 4159, 16)), --  4159 / 0x103f
    4690 => std_logic_vector(to_unsigned( 1037, 16)), --  1037 / 0x040d -- last item of row
    4691 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4692 => std_logic_vector(to_unsigned( 2916, 16)), --  2916 / 0x0b64
    4693 => std_logic_vector(to_unsigned( 2362, 16)), --  2362 / 0x093a -- last item of row
    4694 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4695 => std_logic_vector(to_unsigned(  395, 16)), --   395 / 0x018b
    4696 => std_logic_vector(to_unsigned( 1226, 16)), --  1226 / 0x04ca -- last item of row
    4697 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4698 => std_logic_vector(to_unsigned( 6911, 16)), --  6911 / 0x1aff
    4699 => std_logic_vector(to_unsigned( 4548, 16)), --  4548 / 0x11c4 -- last item of row
    4700 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4701 => std_logic_vector(to_unsigned( 4618, 16)), --  4618 / 0x120a
    4702 => std_logic_vector(to_unsigned( 2241, 16)), --  2241 / 0x08c1 -- last item of row
    4703 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4704 => std_logic_vector(to_unsigned( 4120, 16)), --  4120 / 0x1018
    4705 => std_logic_vector(to_unsigned( 4280, 16)), --  4280 / 0x10b8 -- last item of row
    4706 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4707 => std_logic_vector(to_unsigned( 5825, 16)), --  5825 / 0x16c1
    4708 => std_logic_vector(to_unsigned(  474, 16)), --   474 / 0x01da -- last item of row
    4709 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4710 => std_logic_vector(to_unsigned( 2154, 16)), --  2154 / 0x086a
    4711 => std_logic_vector(to_unsigned( 5558, 16)), --  5558 / 0x15b6 -- last item of row
    4712 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4713 => std_logic_vector(to_unsigned( 3793, 16)), --  3793 / 0x0ed1
    4714 => std_logic_vector(to_unsigned( 5471, 16)), --  5471 / 0x155f -- last item of row
    4715 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4716 => std_logic_vector(to_unsigned( 5707, 16)), --  5707 / 0x164b
    4717 => std_logic_vector(to_unsigned( 1595, 16)), --  1595 / 0x063b -- last item of row
    4718 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4719 => std_logic_vector(to_unsigned( 1403, 16)), --  1403 / 0x057b
    4720 => std_logic_vector(to_unsigned(  325, 16)), --   325 / 0x0145 -- last item of row
    4721 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4722 => std_logic_vector(to_unsigned( 6601, 16)), --  6601 / 0x19c9
    4723 => std_logic_vector(to_unsigned( 5183, 16)), --  5183 / 0x143f -- last item of row
    4724 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4725 => std_logic_vector(to_unsigned( 6369, 16)), --  6369 / 0x18e1
    4726 => std_logic_vector(to_unsigned( 4569, 16)), --  4569 / 0x11d9 -- last item of row
    4727 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4728 => std_logic_vector(to_unsigned( 4846, 16)), --  4846 / 0x12ee
    4729 => std_logic_vector(to_unsigned(  896, 16)), --   896 / 0x0380 -- last item of row
    4730 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4731 => std_logic_vector(to_unsigned( 7092, 16)), --  7092 / 0x1bb4
    4732 => std_logic_vector(to_unsigned( 6184, 16)), --  6184 / 0x1828 -- last item of row
    4733 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4734 => std_logic_vector(to_unsigned( 6764, 16)), --  6764 / 0x1a6c
    4735 => std_logic_vector(to_unsigned( 7127, 16)), --  7127 / 0x1bd7 -- last item of row
    4736 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4737 => std_logic_vector(to_unsigned( 6358, 16)), --  6358 / 0x18d6
    4738 => std_logic_vector(to_unsigned( 1951, 16)), --  1951 / 0x079f -- last item of row
    4739 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4740 => std_logic_vector(to_unsigned( 3117, 16)), --  3117 / 0x0c2d
    4741 => std_logic_vector(to_unsigned( 6960, 16)), --  6960 / 0x1b30 -- last item of row
    4742 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4743 => std_logic_vector(to_unsigned( 2710, 16)), --  2710 / 0x0a96
    4744 => std_logic_vector(to_unsigned( 7062, 16)), --  7062 / 0x1b96 -- last item of row
    4745 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4746 => std_logic_vector(to_unsigned( 1133, 16)), --  1133 / 0x046d
    4747 => std_logic_vector(to_unsigned( 3604, 16)), --  3604 / 0x0e14 -- last item of row
    4748 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4749 => std_logic_vector(to_unsigned( 3694, 16)), --  3694 / 0x0e6e
    4750 => std_logic_vector(to_unsigned(  657, 16)), --   657 / 0x0291 -- last item of row
    4751 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4752 => std_logic_vector(to_unsigned( 1355, 16)), --  1355 / 0x054b
    4753 => std_logic_vector(to_unsigned(  110, 16)), --   110 / 0x006e -- last item of row
    4754 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4755 => std_logic_vector(to_unsigned( 3329, 16)), --  3329 / 0x0d01
    4756 => std_logic_vector(to_unsigned( 6736, 16)), --  6736 / 0x1a50 -- last item of row
    4757 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4758 => std_logic_vector(to_unsigned( 2505, 16)), --  2505 / 0x09c9
    4759 => std_logic_vector(to_unsigned( 3407, 16)), --  3407 / 0x0d4f -- last item of row
    4760 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4761 => std_logic_vector(to_unsigned( 2462, 16)), --  2462 / 0x099e
    4762 => std_logic_vector(to_unsigned( 4806, 16)), --  4806 / 0x12c6 -- last item of row
    4763 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4764 => std_logic_vector(to_unsigned( 4216, 16)), --  4216 / 0x1078
    4765 => std_logic_vector(to_unsigned(  214, 16)), --   214 / 0x00d6 -- last item of row
    4766 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4767 => std_logic_vector(to_unsigned( 5348, 16)), --  5348 / 0x14e4
    4768 => std_logic_vector(to_unsigned( 5619, 16)), --  5619 / 0x15f3 -- last item of row
    4769 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4770 => std_logic_vector(to_unsigned( 6627, 16)), --  6627 / 0x19e3
    4771 => std_logic_vector(to_unsigned( 6243, 16)), --  6243 / 0x1863 -- last item of row
    4772 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4773 => std_logic_vector(to_unsigned( 2644, 16)), --  2644 / 0x0a54
    4774 => std_logic_vector(to_unsigned( 5073, 16)), --  5073 / 0x13d1 -- last item of row
    4775 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4776 => std_logic_vector(to_unsigned( 4212, 16)), --  4212 / 0x1074
    4777 => std_logic_vector(to_unsigned( 5088, 16)), --  5088 / 0x13e0 -- last item of row
    4778 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4779 => std_logic_vector(to_unsigned( 3463, 16)), --  3463 / 0x0d87
    4780 => std_logic_vector(to_unsigned( 3889, 16)), --  3889 / 0x0f31 -- last item of row
    4781 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4782 => std_logic_vector(to_unsigned( 5306, 16)), --  5306 / 0x14ba
    4783 => std_logic_vector(to_unsigned(  478, 16)), --   478 / 0x01de -- last item of row
    4784 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4785 => std_logic_vector(to_unsigned( 4320, 16)), --  4320 / 0x10e0
    4786 => std_logic_vector(to_unsigned( 6121, 16)), --  6121 / 0x17e9 -- last item of row
    4787 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4788 => std_logic_vector(to_unsigned( 3961, 16)), --  3961 / 0x0f79
    4789 => std_logic_vector(to_unsigned( 1125, 16)), --  1125 / 0x0465 -- last item of row
    4790 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4791 => std_logic_vector(to_unsigned( 5699, 16)), --  5699 / 0x1643
    4792 => std_logic_vector(to_unsigned( 1195, 16)), --  1195 / 0x04ab -- last item of row
    4793 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4794 => std_logic_vector(to_unsigned( 6511, 16)), --  6511 / 0x196f
    4795 => std_logic_vector(to_unsigned(  792, 16)), --   792 / 0x0318 -- last item of row
    4796 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4797 => std_logic_vector(to_unsigned( 3934, 16)), --  3934 / 0x0f5e
    4798 => std_logic_vector(to_unsigned( 2778, 16)), --  2778 / 0x0ada -- last item of row
    4799 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4800 => std_logic_vector(to_unsigned( 3238, 16)), --  3238 / 0x0ca6
    4801 => std_logic_vector(to_unsigned( 6587, 16)), --  6587 / 0x19bb -- last item of row
    4802 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4803 => std_logic_vector(to_unsigned( 1111, 16)), --  1111 / 0x0457
    4804 => std_logic_vector(to_unsigned( 6596, 16)), --  6596 / 0x19c4 -- last item of row
    4805 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4806 => std_logic_vector(to_unsigned( 1457, 16)), --  1457 / 0x05b1
    4807 => std_logic_vector(to_unsigned( 6226, 16)), --  6226 / 0x1852 -- last item of row
    4808 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4809 => std_logic_vector(to_unsigned( 1446, 16)), --  1446 / 0x05a6
    4810 => std_logic_vector(to_unsigned( 3885, 16)), --  3885 / 0x0f2d -- last item of row
    4811 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4812 => std_logic_vector(to_unsigned( 3907, 16)), --  3907 / 0x0f43
    4813 => std_logic_vector(to_unsigned( 4043, 16)), --  4043 / 0x0fcb -- last item of row
    4814 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4815 => std_logic_vector(to_unsigned( 6839, 16)), --  6839 / 0x1ab7
    4816 => std_logic_vector(to_unsigned( 2873, 16)), --  2873 / 0x0b39 -- last item of row
    4817 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4818 => std_logic_vector(to_unsigned( 1733, 16)), --  1733 / 0x06c5
    4819 => std_logic_vector(to_unsigned( 5615, 16)), --  5615 / 0x15ef -- last item of row
    4820 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4821 => std_logic_vector(to_unsigned( 5202, 16)), --  5202 / 0x1452
    4822 => std_logic_vector(to_unsigned( 4269, 16)), --  4269 / 0x10ad -- last item of row
    4823 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4824 => std_logic_vector(to_unsigned( 3024, 16)), --  3024 / 0x0bd0
    4825 => std_logic_vector(to_unsigned( 4722, 16)), --  4722 / 0x1272 -- last item of row
    4826 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4827 => std_logic_vector(to_unsigned( 5445, 16)), --  5445 / 0x1545
    4828 => std_logic_vector(to_unsigned( 6372, 16)), --  6372 / 0x18e4 -- last item of row
    4829 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4830 => std_logic_vector(to_unsigned(  370, 16)), --   370 / 0x0172
    4831 => std_logic_vector(to_unsigned( 1828, 16)), --  1828 / 0x0724 -- last item of row
    4832 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4833 => std_logic_vector(to_unsigned( 4695, 16)), --  4695 / 0x1257
    4834 => std_logic_vector(to_unsigned( 1600, 16)), --  1600 / 0x0640 -- last item of row
    4835 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4836 => std_logic_vector(to_unsigned(  680, 16)), --   680 / 0x02a8
    4837 => std_logic_vector(to_unsigned( 2074, 16)), --  2074 / 0x081a -- last item of row
    4838 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4839 => std_logic_vector(to_unsigned( 1801, 16)), --  1801 / 0x0709
    4840 => std_logic_vector(to_unsigned( 6690, 16)), --  6690 / 0x1a22 -- last item of row
    4841 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4842 => std_logic_vector(to_unsigned( 2669, 16)), --  2669 / 0x0a6d
    4843 => std_logic_vector(to_unsigned( 1377, 16)), --  1377 / 0x0561 -- last item of row
    4844 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4845 => std_logic_vector(to_unsigned( 2463, 16)), --  2463 / 0x099f
    4846 => std_logic_vector(to_unsigned( 1681, 16)), --  1681 / 0x0691 -- last item of row
    4847 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4848 => std_logic_vector(to_unsigned( 5972, 16)), --  5972 / 0x1754
    4849 => std_logic_vector(to_unsigned( 5171, 16)), --  5171 / 0x1433 -- last item of row
    4850 => std_logic_vector(to_unsigned(   18, 16)), --    18 / 0x0012
    4851 => std_logic_vector(to_unsigned( 5728, 16)), --  5728 / 0x1660
    4852 => std_logic_vector(to_unsigned( 4284, 16)), --  4284 / 0x10bc -- last item of row
    4853 => std_logic_vector(to_unsigned(   19, 16)), --    19 / 0x0013
    4854 => std_logic_vector(to_unsigned( 1696, 16)), --  1696 / 0x06a0
    4855 => std_logic_vector(to_unsigned( 1459, 16)), --  1459 / 0x05b3 -- last item of row
    -- Table for fecframe_normal, C9_10
    4856 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4857 => std_logic_vector(to_unsigned( 5611, 16)), --  5611 / 0x15eb
    4858 => std_logic_vector(to_unsigned( 2563, 16)), --  2563 / 0x0a03
    4859 => std_logic_vector(to_unsigned( 2900, 16)), --  2900 / 0x0b54 -- last item of row
    4860 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4861 => std_logic_vector(to_unsigned( 5220, 16)), --  5220 / 0x1464
    4862 => std_logic_vector(to_unsigned( 3143, 16)), --  3143 / 0x0c47
    4863 => std_logic_vector(to_unsigned( 4813, 16)), --  4813 / 0x12cd -- last item of row
    4864 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4865 => std_logic_vector(to_unsigned( 2481, 16)), --  2481 / 0x09b1
    4866 => std_logic_vector(to_unsigned(  834, 16)), --   834 / 0x0342
    4867 => std_logic_vector(to_unsigned(   81, 16)), --    81 / 0x0051 -- last item of row
    4868 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4869 => std_logic_vector(to_unsigned( 6265, 16)), --  6265 / 0x1879
    4870 => std_logic_vector(to_unsigned( 4064, 16)), --  4064 / 0x0fe0
    4871 => std_logic_vector(to_unsigned( 4265, 16)), --  4265 / 0x10a9 -- last item of row
    4872 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4873 => std_logic_vector(to_unsigned( 1055, 16)), --  1055 / 0x041f
    4874 => std_logic_vector(to_unsigned( 2914, 16)), --  2914 / 0x0b62
    4875 => std_logic_vector(to_unsigned( 5638, 16)), --  5638 / 0x1606 -- last item of row
    4876 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4877 => std_logic_vector(to_unsigned( 1734, 16)), --  1734 / 0x06c6
    4878 => std_logic_vector(to_unsigned( 2182, 16)), --  2182 / 0x0886
    4879 => std_logic_vector(to_unsigned( 3315, 16)), --  3315 / 0x0cf3 -- last item of row
    4880 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4881 => std_logic_vector(to_unsigned( 3342, 16)), --  3342 / 0x0d0e
    4882 => std_logic_vector(to_unsigned( 5678, 16)), --  5678 / 0x162e
    4883 => std_logic_vector(to_unsigned( 2246, 16)), --  2246 / 0x08c6 -- last item of row
    4884 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4885 => std_logic_vector(to_unsigned( 2185, 16)), --  2185 / 0x0889
    4886 => std_logic_vector(to_unsigned(  552, 16)), --   552 / 0x0228
    4887 => std_logic_vector(to_unsigned( 3385, 16)), --  3385 / 0x0d39 -- last item of row
    4888 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4889 => std_logic_vector(to_unsigned( 2615, 16)), --  2615 / 0x0a37
    4890 => std_logic_vector(to_unsigned(  236, 16)), --   236 / 0x00ec
    4891 => std_logic_vector(to_unsigned( 5334, 16)), --  5334 / 0x14d6 -- last item of row
    4892 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4893 => std_logic_vector(to_unsigned( 1546, 16)), --  1546 / 0x060a
    4894 => std_logic_vector(to_unsigned( 1755, 16)), --  1755 / 0x06db
    4895 => std_logic_vector(to_unsigned( 3846, 16)), --  3846 / 0x0f06 -- last item of row
    4896 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4897 => std_logic_vector(to_unsigned( 4154, 16)), --  4154 / 0x103a
    4898 => std_logic_vector(to_unsigned( 5561, 16)), --  5561 / 0x15b9
    4899 => std_logic_vector(to_unsigned( 3142, 16)), --  3142 / 0x0c46 -- last item of row
    4900 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4901 => std_logic_vector(to_unsigned( 4382, 16)), --  4382 / 0x111e
    4902 => std_logic_vector(to_unsigned( 2957, 16)), --  2957 / 0x0b8d
    4903 => std_logic_vector(to_unsigned( 5400, 16)), --  5400 / 0x1518 -- last item of row
    4904 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4905 => std_logic_vector(to_unsigned( 1209, 16)), --  1209 / 0x04b9
    4906 => std_logic_vector(to_unsigned( 5329, 16)), --  5329 / 0x14d1
    4907 => std_logic_vector(to_unsigned( 3179, 16)), --  3179 / 0x0c6b -- last item of row
    4908 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4909 => std_logic_vector(to_unsigned( 1421, 16)), --  1421 / 0x058d
    4910 => std_logic_vector(to_unsigned( 3528, 16)), --  3528 / 0x0dc8
    4911 => std_logic_vector(to_unsigned( 6063, 16)), --  6063 / 0x17af -- last item of row
    4912 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4913 => std_logic_vector(to_unsigned( 1480, 16)), --  1480 / 0x05c8
    4914 => std_logic_vector(to_unsigned( 1072, 16)), --  1072 / 0x0430
    4915 => std_logic_vector(to_unsigned( 5398, 16)), --  5398 / 0x1516 -- last item of row
    4916 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4917 => std_logic_vector(to_unsigned( 3843, 16)), --  3843 / 0x0f03
    4918 => std_logic_vector(to_unsigned( 1777, 16)), --  1777 / 0x06f1
    4919 => std_logic_vector(to_unsigned( 4369, 16)), --  4369 / 0x1111 -- last item of row
    4920 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4921 => std_logic_vector(to_unsigned( 1334, 16)), --  1334 / 0x0536
    4922 => std_logic_vector(to_unsigned( 2145, 16)), --  2145 / 0x0861
    4923 => std_logic_vector(to_unsigned( 4163, 16)), --  4163 / 0x1043 -- last item of row
    4924 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4925 => std_logic_vector(to_unsigned( 2368, 16)), --  2368 / 0x0940
    4926 => std_logic_vector(to_unsigned( 5055, 16)), --  5055 / 0x13bf
    4927 => std_logic_vector(to_unsigned(  260, 16)), --   260 / 0x0104 -- last item of row
    4928 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4929 => std_logic_vector(to_unsigned( 6118, 16)), --  6118 / 0x17e6
    4930 => std_logic_vector(to_unsigned( 5405, 16)), --  5405 / 0x151d -- last item of row
    4931 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4932 => std_logic_vector(to_unsigned( 2994, 16)), --  2994 / 0x0bb2
    4933 => std_logic_vector(to_unsigned( 4370, 16)), --  4370 / 0x1112 -- last item of row
    4934 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4935 => std_logic_vector(to_unsigned( 3405, 16)), --  3405 / 0x0d4d
    4936 => std_logic_vector(to_unsigned( 1669, 16)), --  1669 / 0x0685 -- last item of row
    4937 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4938 => std_logic_vector(to_unsigned( 4640, 16)), --  4640 / 0x1220
    4939 => std_logic_vector(to_unsigned( 5550, 16)), --  5550 / 0x15ae -- last item of row
    4940 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4941 => std_logic_vector(to_unsigned( 1354, 16)), --  1354 / 0x054a
    4942 => std_logic_vector(to_unsigned( 3921, 16)), --  3921 / 0x0f51 -- last item of row
    4943 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4944 => std_logic_vector(to_unsigned(  117, 16)), --   117 / 0x0075
    4945 => std_logic_vector(to_unsigned( 1713, 16)), --  1713 / 0x06b1 -- last item of row
    4946 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    4947 => std_logic_vector(to_unsigned( 5425, 16)), --  5425 / 0x1531
    4948 => std_logic_vector(to_unsigned( 2866, 16)), --  2866 / 0x0b32 -- last item of row
    4949 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    4950 => std_logic_vector(to_unsigned( 6047, 16)), --  6047 / 0x179f
    4951 => std_logic_vector(to_unsigned(  683, 16)), --   683 / 0x02ab -- last item of row
    4952 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    4953 => std_logic_vector(to_unsigned( 5616, 16)), --  5616 / 0x15f0
    4954 => std_logic_vector(to_unsigned( 2582, 16)), --  2582 / 0x0a16 -- last item of row
    4955 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    4956 => std_logic_vector(to_unsigned( 2108, 16)), --  2108 / 0x083c
    4957 => std_logic_vector(to_unsigned( 1179, 16)), --  1179 / 0x049b -- last item of row
    4958 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    4959 => std_logic_vector(to_unsigned(  933, 16)), --   933 / 0x03a5
    4960 => std_logic_vector(to_unsigned( 4921, 16)), --  4921 / 0x1339 -- last item of row
    4961 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    4962 => std_logic_vector(to_unsigned( 5953, 16)), --  5953 / 0x1741
    4963 => std_logic_vector(to_unsigned( 2261, 16)), --  2261 / 0x08d5 -- last item of row
    4964 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    4965 => std_logic_vector(to_unsigned( 1430, 16)), --  1430 / 0x0596
    4966 => std_logic_vector(to_unsigned( 4699, 16)), --  4699 / 0x125b -- last item of row
    4967 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    4968 => std_logic_vector(to_unsigned( 5905, 16)), --  5905 / 0x1711
    4969 => std_logic_vector(to_unsigned(  480, 16)), --   480 / 0x01e0 -- last item of row
    4970 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    4971 => std_logic_vector(to_unsigned( 4289, 16)), --  4289 / 0x10c1
    4972 => std_logic_vector(to_unsigned( 1846, 16)), --  1846 / 0x0736 -- last item of row
    4973 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    4974 => std_logic_vector(to_unsigned( 5374, 16)), --  5374 / 0x14fe
    4975 => std_logic_vector(to_unsigned( 6208, 16)), --  6208 / 0x1840 -- last item of row
    4976 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    4977 => std_logic_vector(to_unsigned( 1775, 16)), --  1775 / 0x06ef
    4978 => std_logic_vector(to_unsigned( 3476, 16)), --  3476 / 0x0d94 -- last item of row
    4979 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    4980 => std_logic_vector(to_unsigned( 3216, 16)), --  3216 / 0x0c90
    4981 => std_logic_vector(to_unsigned( 2178, 16)), --  2178 / 0x0882 -- last item of row
    4982 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    4983 => std_logic_vector(to_unsigned( 4165, 16)), --  4165 / 0x1045
    4984 => std_logic_vector(to_unsigned(  884, 16)), --   884 / 0x0374 -- last item of row
    4985 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    4986 => std_logic_vector(to_unsigned( 2896, 16)), --  2896 / 0x0b50
    4987 => std_logic_vector(to_unsigned( 3744, 16)), --  3744 / 0x0ea0 -- last item of row
    4988 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    4989 => std_logic_vector(to_unsigned(  874, 16)), --   874 / 0x036a
    4990 => std_logic_vector(to_unsigned( 2801, 16)), --  2801 / 0x0af1 -- last item of row
    4991 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    4992 => std_logic_vector(to_unsigned( 3423, 16)), --  3423 / 0x0d5f
    4993 => std_logic_vector(to_unsigned( 5579, 16)), --  5579 / 0x15cb -- last item of row
    4994 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    4995 => std_logic_vector(to_unsigned( 3404, 16)), --  3404 / 0x0d4c
    4996 => std_logic_vector(to_unsigned( 3552, 16)), --  3552 / 0x0de0 -- last item of row
    4997 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    4998 => std_logic_vector(to_unsigned( 2876, 16)), --  2876 / 0x0b3c
    4999 => std_logic_vector(to_unsigned( 5515, 16)), --  5515 / 0x158b -- last item of row
    5000 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5001 => std_logic_vector(to_unsigned(  516, 16)), --   516 / 0x0204
    5002 => std_logic_vector(to_unsigned( 1719, 16)), --  1719 / 0x06b7 -- last item of row
    5003 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5004 => std_logic_vector(to_unsigned(  765, 16)), --   765 / 0x02fd
    5005 => std_logic_vector(to_unsigned( 3631, 16)), --  3631 / 0x0e2f -- last item of row
    5006 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5007 => std_logic_vector(to_unsigned( 5059, 16)), --  5059 / 0x13c3
    5008 => std_logic_vector(to_unsigned( 1441, 16)), --  1441 / 0x05a1 -- last item of row
    5009 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5010 => std_logic_vector(to_unsigned( 5629, 16)), --  5629 / 0x15fd
    5011 => std_logic_vector(to_unsigned(  598, 16)), --   598 / 0x0256 -- last item of row
    5012 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5013 => std_logic_vector(to_unsigned( 5405, 16)), --  5405 / 0x151d
    5014 => std_logic_vector(to_unsigned(  473, 16)), --   473 / 0x01d9 -- last item of row
    5015 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5016 => std_logic_vector(to_unsigned( 4724, 16)), --  4724 / 0x1274
    5017 => std_logic_vector(to_unsigned( 5210, 16)), --  5210 / 0x145a -- last item of row
    5018 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5019 => std_logic_vector(to_unsigned(  155, 16)), --   155 / 0x009b
    5020 => std_logic_vector(to_unsigned( 1832, 16)), --  1832 / 0x0728 -- last item of row
    5021 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5022 => std_logic_vector(to_unsigned( 1689, 16)), --  1689 / 0x0699
    5023 => std_logic_vector(to_unsigned( 2229, 16)), --  2229 / 0x08b5 -- last item of row
    5024 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5025 => std_logic_vector(to_unsigned(  449, 16)), --   449 / 0x01c1
    5026 => std_logic_vector(to_unsigned( 1164, 16)), --  1164 / 0x048c -- last item of row
    5027 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5028 => std_logic_vector(to_unsigned( 2308, 16)), --  2308 / 0x0904
    5029 => std_logic_vector(to_unsigned( 3088, 16)), --  3088 / 0x0c10 -- last item of row
    5030 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5031 => std_logic_vector(to_unsigned( 1122, 16)), --  1122 / 0x0462
    5032 => std_logic_vector(to_unsigned(  669, 16)), --   669 / 0x029d -- last item of row
    5033 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5034 => std_logic_vector(to_unsigned( 2268, 16)), --  2268 / 0x08dc
    5035 => std_logic_vector(to_unsigned( 5758, 16)), --  5758 / 0x167e -- last item of row
    5036 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5037 => std_logic_vector(to_unsigned( 5878, 16)), --  5878 / 0x16f6
    5038 => std_logic_vector(to_unsigned( 2609, 16)), --  2609 / 0x0a31 -- last item of row
    5039 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5040 => std_logic_vector(to_unsigned(  782, 16)), --   782 / 0x030e
    5041 => std_logic_vector(to_unsigned( 3359, 16)), --  3359 / 0x0d1f -- last item of row
    5042 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5043 => std_logic_vector(to_unsigned( 1231, 16)), --  1231 / 0x04cf
    5044 => std_logic_vector(to_unsigned( 4231, 16)), --  4231 / 0x1087 -- last item of row
    5045 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5046 => std_logic_vector(to_unsigned( 4225, 16)), --  4225 / 0x1081
    5047 => std_logic_vector(to_unsigned( 2052, 16)), --  2052 / 0x0804 -- last item of row
    5048 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5049 => std_logic_vector(to_unsigned( 4286, 16)), --  4286 / 0x10be
    5050 => std_logic_vector(to_unsigned( 3517, 16)), --  3517 / 0x0dbd -- last item of row
    5051 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5052 => std_logic_vector(to_unsigned( 5531, 16)), --  5531 / 0x159b
    5053 => std_logic_vector(to_unsigned( 3184, 16)), --  3184 / 0x0c70 -- last item of row
    5054 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5055 => std_logic_vector(to_unsigned( 1935, 16)), --  1935 / 0x078f
    5056 => std_logic_vector(to_unsigned( 4560, 16)), --  4560 / 0x11d0 -- last item of row
    5057 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5058 => std_logic_vector(to_unsigned( 1174, 16)), --  1174 / 0x0496
    5059 => std_logic_vector(to_unsigned(  131, 16)), --   131 / 0x0083 -- last item of row
    5060 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5061 => std_logic_vector(to_unsigned( 3115, 16)), --  3115 / 0x0c2b
    5062 => std_logic_vector(to_unsigned(  956, 16)), --   956 / 0x03bc -- last item of row
    5063 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5064 => std_logic_vector(to_unsigned( 3129, 16)), --  3129 / 0x0c39
    5065 => std_logic_vector(to_unsigned( 1088, 16)), --  1088 / 0x0440 -- last item of row
    5066 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5067 => std_logic_vector(to_unsigned( 5238, 16)), --  5238 / 0x1476
    5068 => std_logic_vector(to_unsigned( 4440, 16)), --  4440 / 0x1158 -- last item of row
    5069 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5070 => std_logic_vector(to_unsigned( 5722, 16)), --  5722 / 0x165a
    5071 => std_logic_vector(to_unsigned( 4280, 16)), --  4280 / 0x10b8 -- last item of row
    5072 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5073 => std_logic_vector(to_unsigned( 3540, 16)), --  3540 / 0x0dd4
    5074 => std_logic_vector(to_unsigned(  375, 16)), --   375 / 0x0177 -- last item of row
    5075 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5076 => std_logic_vector(to_unsigned(  191, 16)), --   191 / 0x00bf
    5077 => std_logic_vector(to_unsigned( 2782, 16)), --  2782 / 0x0ade -- last item of row
    5078 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5079 => std_logic_vector(to_unsigned(  906, 16)), --   906 / 0x038a
    5080 => std_logic_vector(to_unsigned( 4432, 16)), --  4432 / 0x1150 -- last item of row
    5081 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5082 => std_logic_vector(to_unsigned( 3225, 16)), --  3225 / 0x0c99
    5083 => std_logic_vector(to_unsigned( 1111, 16)), --  1111 / 0x0457 -- last item of row
    5084 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5085 => std_logic_vector(to_unsigned( 6296, 16)), --  6296 / 0x1898
    5086 => std_logic_vector(to_unsigned( 2583, 16)), --  2583 / 0x0a17 -- last item of row
    5087 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5088 => std_logic_vector(to_unsigned( 1457, 16)), --  1457 / 0x05b1
    5089 => std_logic_vector(to_unsigned(  903, 16)), --   903 / 0x0387 -- last item of row
    5090 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5091 => std_logic_vector(to_unsigned(  855, 16)), --   855 / 0x0357
    5092 => std_logic_vector(to_unsigned( 4475, 16)), --  4475 / 0x117b -- last item of row
    5093 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5094 => std_logic_vector(to_unsigned( 4097, 16)), --  4097 / 0x1001
    5095 => std_logic_vector(to_unsigned( 3970, 16)), --  3970 / 0x0f82 -- last item of row
    5096 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5097 => std_logic_vector(to_unsigned( 4433, 16)), --  4433 / 0x1151
    5098 => std_logic_vector(to_unsigned( 4361, 16)), --  4361 / 0x1109 -- last item of row
    5099 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5100 => std_logic_vector(to_unsigned( 5198, 16)), --  5198 / 0x144e
    5101 => std_logic_vector(to_unsigned(  541, 16)), --   541 / 0x021d -- last item of row
    5102 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5103 => std_logic_vector(to_unsigned( 1146, 16)), --  1146 / 0x047a
    5104 => std_logic_vector(to_unsigned( 4426, 16)), --  4426 / 0x114a -- last item of row
    5105 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5106 => std_logic_vector(to_unsigned( 3202, 16)), --  3202 / 0x0c82
    5107 => std_logic_vector(to_unsigned( 2902, 16)), --  2902 / 0x0b56 -- last item of row
    5108 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5109 => std_logic_vector(to_unsigned( 2724, 16)), --  2724 / 0x0aa4
    5110 => std_logic_vector(to_unsigned(  525, 16)), --   525 / 0x020d -- last item of row
    5111 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5112 => std_logic_vector(to_unsigned( 1083, 16)), --  1083 / 0x043b
    5113 => std_logic_vector(to_unsigned( 4124, 16)), --  4124 / 0x101c -- last item of row
    5114 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5115 => std_logic_vector(to_unsigned( 2326, 16)), --  2326 / 0x0916
    5116 => std_logic_vector(to_unsigned( 6003, 16)), --  6003 / 0x1773 -- last item of row
    5117 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5118 => std_logic_vector(to_unsigned( 5605, 16)), --  5605 / 0x15e5
    5119 => std_logic_vector(to_unsigned( 5990, 16)), --  5990 / 0x1766 -- last item of row
    5120 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5121 => std_logic_vector(to_unsigned( 4376, 16)), --  4376 / 0x1118
    5122 => std_logic_vector(to_unsigned( 1579, 16)), --  1579 / 0x062b -- last item of row
    5123 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5124 => std_logic_vector(to_unsigned( 4407, 16)), --  4407 / 0x1137
    5125 => std_logic_vector(to_unsigned(  984, 16)), --   984 / 0x03d8 -- last item of row
    5126 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5127 => std_logic_vector(to_unsigned( 1332, 16)), --  1332 / 0x0534
    5128 => std_logic_vector(to_unsigned( 6163, 16)), --  6163 / 0x1813 -- last item of row
    5129 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5130 => std_logic_vector(to_unsigned( 5359, 16)), --  5359 / 0x14ef
    5131 => std_logic_vector(to_unsigned( 3975, 16)), --  3975 / 0x0f87 -- last item of row
    5132 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5133 => std_logic_vector(to_unsigned( 1907, 16)), --  1907 / 0x0773
    5134 => std_logic_vector(to_unsigned( 1854, 16)), --  1854 / 0x073e -- last item of row
    5135 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5136 => std_logic_vector(to_unsigned( 3601, 16)), --  3601 / 0x0e11
    5137 => std_logic_vector(to_unsigned( 5748, 16)), --  5748 / 0x1674 -- last item of row
    5138 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5139 => std_logic_vector(to_unsigned( 6056, 16)), --  6056 / 0x17a8
    5140 => std_logic_vector(to_unsigned( 3266, 16)), --  3266 / 0x0cc2 -- last item of row
    5141 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5142 => std_logic_vector(to_unsigned( 3322, 16)), --  3322 / 0x0cfa
    5143 => std_logic_vector(to_unsigned( 4085, 16)), --  4085 / 0x0ff5 -- last item of row
    5144 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5145 => std_logic_vector(to_unsigned( 1768, 16)), --  1768 / 0x06e8
    5146 => std_logic_vector(to_unsigned( 3244, 16)), --  3244 / 0x0cac -- last item of row
    5147 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5148 => std_logic_vector(to_unsigned( 2149, 16)), --  2149 / 0x0865
    5149 => std_logic_vector(to_unsigned(  144, 16)), --   144 / 0x0090 -- last item of row
    5150 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5151 => std_logic_vector(to_unsigned( 1589, 16)), --  1589 / 0x0635
    5152 => std_logic_vector(to_unsigned( 4291, 16)), --  4291 / 0x10c3 -- last item of row
    5153 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5154 => std_logic_vector(to_unsigned( 5154, 16)), --  5154 / 0x1422
    5155 => std_logic_vector(to_unsigned( 1252, 16)), --  1252 / 0x04e4 -- last item of row
    5156 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5157 => std_logic_vector(to_unsigned( 1855, 16)), --  1855 / 0x073f
    5158 => std_logic_vector(to_unsigned( 5939, 16)), --  5939 / 0x1733 -- last item of row
    5159 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5160 => std_logic_vector(to_unsigned( 4820, 16)), --  4820 / 0x12d4
    5161 => std_logic_vector(to_unsigned( 2706, 16)), --  2706 / 0x0a92 -- last item of row
    5162 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5163 => std_logic_vector(to_unsigned( 1475, 16)), --  1475 / 0x05c3
    5164 => std_logic_vector(to_unsigned( 3360, 16)), --  3360 / 0x0d20 -- last item of row
    5165 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5166 => std_logic_vector(to_unsigned( 4266, 16)), --  4266 / 0x10aa
    5167 => std_logic_vector(to_unsigned(  693, 16)), --   693 / 0x02b5 -- last item of row
    5168 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5169 => std_logic_vector(to_unsigned( 4156, 16)), --  4156 / 0x103c
    5170 => std_logic_vector(to_unsigned( 2018, 16)), --  2018 / 0x07e2 -- last item of row
    5171 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5172 => std_logic_vector(to_unsigned( 2103, 16)), --  2103 / 0x0837
    5173 => std_logic_vector(to_unsigned(  752, 16)), --   752 / 0x02f0 -- last item of row
    5174 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5175 => std_logic_vector(to_unsigned( 3710, 16)), --  3710 / 0x0e7e
    5176 => std_logic_vector(to_unsigned( 3853, 16)), --  3853 / 0x0f0d -- last item of row
    5177 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5178 => std_logic_vector(to_unsigned( 5123, 16)), --  5123 / 0x1403
    5179 => std_logic_vector(to_unsigned(  931, 16)), --   931 / 0x03a3 -- last item of row
    5180 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5181 => std_logic_vector(to_unsigned( 6146, 16)), --  6146 / 0x1802
    5182 => std_logic_vector(to_unsigned( 3323, 16)), --  3323 / 0x0cfb -- last item of row
    5183 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5184 => std_logic_vector(to_unsigned( 1939, 16)), --  1939 / 0x0793
    5185 => std_logic_vector(to_unsigned( 5002, 16)), --  5002 / 0x138a -- last item of row
    5186 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5187 => std_logic_vector(to_unsigned( 5140, 16)), --  5140 / 0x1414
    5188 => std_logic_vector(to_unsigned( 1437, 16)), --  1437 / 0x059d -- last item of row
    5189 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5190 => std_logic_vector(to_unsigned( 1263, 16)), --  1263 / 0x04ef
    5191 => std_logic_vector(to_unsigned(  293, 16)), --   293 / 0x0125 -- last item of row
    5192 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5193 => std_logic_vector(to_unsigned( 5949, 16)), --  5949 / 0x173d
    5194 => std_logic_vector(to_unsigned( 4665, 16)), --  4665 / 0x1239 -- last item of row
    5195 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5196 => std_logic_vector(to_unsigned( 4548, 16)), --  4548 / 0x11c4
    5197 => std_logic_vector(to_unsigned( 6380, 16)), --  6380 / 0x18ec -- last item of row
    5198 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5199 => std_logic_vector(to_unsigned( 3171, 16)), --  3171 / 0x0c63
    5200 => std_logic_vector(to_unsigned( 4690, 16)), --  4690 / 0x1252 -- last item of row
    5201 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5202 => std_logic_vector(to_unsigned( 5204, 16)), --  5204 / 0x1454
    5203 => std_logic_vector(to_unsigned( 2114, 16)), --  2114 / 0x0842 -- last item of row
    5204 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5205 => std_logic_vector(to_unsigned( 6384, 16)), --  6384 / 0x18f0
    5206 => std_logic_vector(to_unsigned( 5565, 16)), --  5565 / 0x15bd -- last item of row
    5207 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5208 => std_logic_vector(to_unsigned( 5722, 16)), --  5722 / 0x165a
    5209 => std_logic_vector(to_unsigned( 1757, 16)), --  1757 / 0x06dd -- last item of row
    5210 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5211 => std_logic_vector(to_unsigned( 2805, 16)), --  2805 / 0x0af5
    5212 => std_logic_vector(to_unsigned( 6264, 16)), --  6264 / 0x1878 -- last item of row
    5213 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5214 => std_logic_vector(to_unsigned( 1202, 16)), --  1202 / 0x04b2
    5215 => std_logic_vector(to_unsigned( 2616, 16)), --  2616 / 0x0a38 -- last item of row
    5216 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5217 => std_logic_vector(to_unsigned( 1018, 16)), --  1018 / 0x03fa
    5218 => std_logic_vector(to_unsigned( 3244, 16)), --  3244 / 0x0cac -- last item of row
    5219 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5220 => std_logic_vector(to_unsigned( 4018, 16)), --  4018 / 0x0fb2
    5221 => std_logic_vector(to_unsigned( 5289, 16)), --  5289 / 0x14a9 -- last item of row
    5222 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5223 => std_logic_vector(to_unsigned( 2257, 16)), --  2257 / 0x08d1
    5224 => std_logic_vector(to_unsigned( 3067, 16)), --  3067 / 0x0bfb -- last item of row
    5225 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5226 => std_logic_vector(to_unsigned( 2483, 16)), --  2483 / 0x09b3
    5227 => std_logic_vector(to_unsigned( 3073, 16)), --  3073 / 0x0c01 -- last item of row
    5228 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5229 => std_logic_vector(to_unsigned( 1196, 16)), --  1196 / 0x04ac
    5230 => std_logic_vector(to_unsigned( 5329, 16)), --  5329 / 0x14d1 -- last item of row
    5231 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5232 => std_logic_vector(to_unsigned(  649, 16)), --   649 / 0x0289
    5233 => std_logic_vector(to_unsigned( 3918, 16)), --  3918 / 0x0f4e -- last item of row
    5234 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5235 => std_logic_vector(to_unsigned( 3791, 16)), --  3791 / 0x0ecf
    5236 => std_logic_vector(to_unsigned( 4581, 16)), --  4581 / 0x11e5 -- last item of row
    5237 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5238 => std_logic_vector(to_unsigned( 5028, 16)), --  5028 / 0x13a4
    5239 => std_logic_vector(to_unsigned( 3803, 16)), --  3803 / 0x0edb -- last item of row
    5240 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5241 => std_logic_vector(to_unsigned( 3119, 16)), --  3119 / 0x0c2f
    5242 => std_logic_vector(to_unsigned( 3506, 16)), --  3506 / 0x0db2 -- last item of row
    5243 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5244 => std_logic_vector(to_unsigned( 4779, 16)), --  4779 / 0x12ab
    5245 => std_logic_vector(to_unsigned(  431, 16)), --   431 / 0x01af -- last item of row
    5246 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5247 => std_logic_vector(to_unsigned( 3888, 16)), --  3888 / 0x0f30
    5248 => std_logic_vector(to_unsigned( 5510, 16)), --  5510 / 0x1586 -- last item of row
    5249 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5250 => std_logic_vector(to_unsigned( 4387, 16)), --  4387 / 0x1123
    5251 => std_logic_vector(to_unsigned( 4084, 16)), --  4084 / 0x0ff4 -- last item of row
    5252 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5253 => std_logic_vector(to_unsigned( 5836, 16)), --  5836 / 0x16cc
    5254 => std_logic_vector(to_unsigned( 1692, 16)), --  1692 / 0x069c -- last item of row
    5255 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5256 => std_logic_vector(to_unsigned( 5126, 16)), --  5126 / 0x1406
    5257 => std_logic_vector(to_unsigned( 1078, 16)), --  1078 / 0x0436 -- last item of row
    5258 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5259 => std_logic_vector(to_unsigned( 5721, 16)), --  5721 / 0x1659
    5260 => std_logic_vector(to_unsigned( 6165, 16)), --  6165 / 0x1815 -- last item of row
    5261 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5262 => std_logic_vector(to_unsigned( 3540, 16)), --  3540 / 0x0dd4
    5263 => std_logic_vector(to_unsigned( 2499, 16)), --  2499 / 0x09c3 -- last item of row
    5264 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5265 => std_logic_vector(to_unsigned( 2225, 16)), --  2225 / 0x08b1
    5266 => std_logic_vector(to_unsigned( 6348, 16)), --  6348 / 0x18cc -- last item of row
    5267 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5268 => std_logic_vector(to_unsigned( 1044, 16)), --  1044 / 0x0414
    5269 => std_logic_vector(to_unsigned( 1484, 16)), --  1484 / 0x05cc -- last item of row
    5270 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5271 => std_logic_vector(to_unsigned( 6323, 16)), --  6323 / 0x18b3
    5272 => std_logic_vector(to_unsigned( 4042, 16)), --  4042 / 0x0fca -- last item of row
    5273 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5274 => std_logic_vector(to_unsigned( 1313, 16)), --  1313 / 0x0521
    5275 => std_logic_vector(to_unsigned( 5603, 16)), --  5603 / 0x15e3 -- last item of row
    5276 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5277 => std_logic_vector(to_unsigned( 1303, 16)), --  1303 / 0x0517
    5278 => std_logic_vector(to_unsigned( 3496, 16)), --  3496 / 0x0da8 -- last item of row
    5279 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5280 => std_logic_vector(to_unsigned( 3516, 16)), --  3516 / 0x0dbc
    5281 => std_logic_vector(to_unsigned( 3639, 16)), --  3639 / 0x0e37 -- last item of row
    5282 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5283 => std_logic_vector(to_unsigned( 5161, 16)), --  5161 / 0x1429
    5284 => std_logic_vector(to_unsigned( 2293, 16)), --  2293 / 0x08f5 -- last item of row
    5285 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5286 => std_logic_vector(to_unsigned( 4682, 16)), --  4682 / 0x124a
    5287 => std_logic_vector(to_unsigned( 3845, 16)), --  3845 / 0x0f05 -- last item of row
    5288 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5289 => std_logic_vector(to_unsigned( 3045, 16)), --  3045 / 0x0be5
    5290 => std_logic_vector(to_unsigned(  643, 16)), --   643 / 0x0283 -- last item of row
    5291 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5292 => std_logic_vector(to_unsigned( 2818, 16)), --  2818 / 0x0b02
    5293 => std_logic_vector(to_unsigned( 2616, 16)), --  2616 / 0x0a38 -- last item of row
    5294 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5295 => std_logic_vector(to_unsigned( 3267, 16)), --  3267 / 0x0cc3
    5296 => std_logic_vector(to_unsigned(  649, 16)), --   649 / 0x0289 -- last item of row
    5297 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5298 => std_logic_vector(to_unsigned( 6236, 16)), --  6236 / 0x185c
    5299 => std_logic_vector(to_unsigned(  593, 16)), --   593 / 0x0251 -- last item of row
    5300 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5301 => std_logic_vector(to_unsigned(  646, 16)), --   646 / 0x0286
    5302 => std_logic_vector(to_unsigned( 2948, 16)), --  2948 / 0x0b84 -- last item of row
    5303 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5304 => std_logic_vector(to_unsigned( 4213, 16)), --  4213 / 0x1075
    5305 => std_logic_vector(to_unsigned( 1442, 16)), --  1442 / 0x05a2 -- last item of row
    5306 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5307 => std_logic_vector(to_unsigned( 5779, 16)), --  5779 / 0x1693
    5308 => std_logic_vector(to_unsigned( 1596, 16)), --  1596 / 0x063c -- last item of row
    5309 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5310 => std_logic_vector(to_unsigned( 2403, 16)), --  2403 / 0x0963
    5311 => std_logic_vector(to_unsigned( 1237, 16)), --  1237 / 0x04d5 -- last item of row
    5312 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5313 => std_logic_vector(to_unsigned( 2217, 16)), --  2217 / 0x08a9
    5314 => std_logic_vector(to_unsigned( 1514, 16)), --  1514 / 0x05ea -- last item of row
    5315 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5316 => std_logic_vector(to_unsigned( 5609, 16)), --  5609 / 0x15e9
    5317 => std_logic_vector(to_unsigned(  716, 16)), --   716 / 0x02cc -- last item of row
    5318 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5319 => std_logic_vector(to_unsigned( 5155, 16)), --  5155 / 0x1423
    5320 => std_logic_vector(to_unsigned( 3858, 16)), --  3858 / 0x0f12 -- last item of row
    5321 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5322 => std_logic_vector(to_unsigned( 1517, 16)), --  1517 / 0x05ed
    5323 => std_logic_vector(to_unsigned( 1312, 16)), --  1312 / 0x0520 -- last item of row
    5324 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5325 => std_logic_vector(to_unsigned( 2554, 16)), --  2554 / 0x09fa
    5326 => std_logic_vector(to_unsigned( 3158, 16)), --  3158 / 0x0c56 -- last item of row
    5327 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5328 => std_logic_vector(to_unsigned( 5280, 16)), --  5280 / 0x14a0
    5329 => std_logic_vector(to_unsigned( 2643, 16)), --  2643 / 0x0a53 -- last item of row
    5330 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5331 => std_logic_vector(to_unsigned( 4990, 16)), --  4990 / 0x137e
    5332 => std_logic_vector(to_unsigned( 1353, 16)), --  1353 / 0x0549 -- last item of row
    5333 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5334 => std_logic_vector(to_unsigned( 5648, 16)), --  5648 / 0x1610
    5335 => std_logic_vector(to_unsigned( 1170, 16)), --  1170 / 0x0492 -- last item of row
    5336 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5337 => std_logic_vector(to_unsigned( 1152, 16)), --  1152 / 0x0480
    5338 => std_logic_vector(to_unsigned( 4366, 16)), --  4366 / 0x110e -- last item of row
    5339 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5340 => std_logic_vector(to_unsigned( 3561, 16)), --  3561 / 0x0de9
    5341 => std_logic_vector(to_unsigned( 5368, 16)), --  5368 / 0x14f8 -- last item of row
    5342 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5343 => std_logic_vector(to_unsigned( 3581, 16)), --  3581 / 0x0dfd
    5344 => std_logic_vector(to_unsigned( 1411, 16)), --  1411 / 0x0583 -- last item of row
    5345 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5346 => std_logic_vector(to_unsigned( 5647, 16)), --  5647 / 0x160f
    5347 => std_logic_vector(to_unsigned( 4661, 16)), --  4661 / 0x1235 -- last item of row
    5348 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5349 => std_logic_vector(to_unsigned( 1542, 16)), --  1542 / 0x0606
    5350 => std_logic_vector(to_unsigned( 5401, 16)), --  5401 / 0x1519 -- last item of row
    5351 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    5352 => std_logic_vector(to_unsigned( 5078, 16)), --  5078 / 0x13d6
    5353 => std_logic_vector(to_unsigned( 2687, 16)), --  2687 / 0x0a7f -- last item of row
    5354 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    5355 => std_logic_vector(to_unsigned(  316, 16)), --   316 / 0x013c
    5356 => std_logic_vector(to_unsigned( 1755, 16)), --  1755 / 0x06db -- last item of row
    5357 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    5358 => std_logic_vector(to_unsigned( 3392, 16)), --  3392 / 0x0d40
    5359 => std_logic_vector(to_unsigned( 1991, 16)), --  1991 / 0x07c7 -- last item of row
    -- Table for fecframe_short, C1_2
    5360 => std_logic_vector(to_unsigned(   20, 16)), --    20 / 0x0014
    5361 => std_logic_vector(to_unsigned(  712, 16)), --   712 / 0x02c8
    5362 => std_logic_vector(to_unsigned( 2386, 16)), --  2386 / 0x0952
    5363 => std_logic_vector(to_unsigned( 6354, 16)), --  6354 / 0x18d2
    5364 => std_logic_vector(to_unsigned( 4061, 16)), --  4061 / 0x0fdd
    5365 => std_logic_vector(to_unsigned( 1062, 16)), --  1062 / 0x0426
    5366 => std_logic_vector(to_unsigned( 5045, 16)), --  5045 / 0x13b5
    5367 => std_logic_vector(to_unsigned( 5158, 16)), --  5158 / 0x1426 -- last item of row
    5368 => std_logic_vector(to_unsigned(   21, 16)), --    21 / 0x0015
    5369 => std_logic_vector(to_unsigned( 2543, 16)), --  2543 / 0x09ef
    5370 => std_logic_vector(to_unsigned( 5748, 16)), --  5748 / 0x1674
    5371 => std_logic_vector(to_unsigned( 4822, 16)), --  4822 / 0x12d6
    5372 => std_logic_vector(to_unsigned( 2348, 16)), --  2348 / 0x092c
    5373 => std_logic_vector(to_unsigned( 3089, 16)), --  3089 / 0x0c11
    5374 => std_logic_vector(to_unsigned( 6328, 16)), --  6328 / 0x18b8
    5375 => std_logic_vector(to_unsigned( 5876, 16)), --  5876 / 0x16f4 -- last item of row
    5376 => std_logic_vector(to_unsigned(   22, 16)), --    22 / 0x0016
    5377 => std_logic_vector(to_unsigned(  926, 16)), --   926 / 0x039e
    5378 => std_logic_vector(to_unsigned( 5701, 16)), --  5701 / 0x1645
    5379 => std_logic_vector(to_unsigned(  269, 16)), --   269 / 0x010d
    5380 => std_logic_vector(to_unsigned( 3693, 16)), --  3693 / 0x0e6d
    5381 => std_logic_vector(to_unsigned( 2438, 16)), --  2438 / 0x0986
    5382 => std_logic_vector(to_unsigned( 3190, 16)), --  3190 / 0x0c76
    5383 => std_logic_vector(to_unsigned( 3507, 16)), --  3507 / 0x0db3 -- last item of row
    5384 => std_logic_vector(to_unsigned(   23, 16)), --    23 / 0x0017
    5385 => std_logic_vector(to_unsigned( 2802, 16)), --  2802 / 0x0af2
    5386 => std_logic_vector(to_unsigned( 4520, 16)), --  4520 / 0x11a8
    5387 => std_logic_vector(to_unsigned( 3577, 16)), --  3577 / 0x0df9
    5388 => std_logic_vector(to_unsigned( 5324, 16)), --  5324 / 0x14cc
    5389 => std_logic_vector(to_unsigned( 1091, 16)), --  1091 / 0x0443
    5390 => std_logic_vector(to_unsigned( 4667, 16)), --  4667 / 0x123b
    5391 => std_logic_vector(to_unsigned( 4449, 16)), --  4449 / 0x1161 -- last item of row
    5392 => std_logic_vector(to_unsigned(   24, 16)), --    24 / 0x0018
    5393 => std_logic_vector(to_unsigned( 5140, 16)), --  5140 / 0x1414
    5394 => std_logic_vector(to_unsigned( 2003, 16)), --  2003 / 0x07d3
    5395 => std_logic_vector(to_unsigned( 1263, 16)), --  1263 / 0x04ef
    5396 => std_logic_vector(to_unsigned( 4742, 16)), --  4742 / 0x1286
    5397 => std_logic_vector(to_unsigned( 6497, 16)), --  6497 / 0x1961
    5398 => std_logic_vector(to_unsigned( 1185, 16)), --  1185 / 0x04a1
    5399 => std_logic_vector(to_unsigned( 6202, 16)), --  6202 / 0x183a -- last item of row
    5400 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5401 => std_logic_vector(to_unsigned( 4046, 16)), --  4046 / 0x0fce
    5402 => std_logic_vector(to_unsigned( 6934, 16)), --  6934 / 0x1b16 -- last item of row
    5403 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5404 => std_logic_vector(to_unsigned( 2855, 16)), --  2855 / 0x0b27
    5405 => std_logic_vector(to_unsigned(   66, 16)), --    66 / 0x0042 -- last item of row
    5406 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5407 => std_logic_vector(to_unsigned( 6694, 16)), --  6694 / 0x1a26
    5408 => std_logic_vector(to_unsigned(  212, 16)), --   212 / 0x00d4 -- last item of row
    5409 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5410 => std_logic_vector(to_unsigned( 3439, 16)), --  3439 / 0x0d6f
    5411 => std_logic_vector(to_unsigned( 1158, 16)), --  1158 / 0x0486 -- last item of row
    5412 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5413 => std_logic_vector(to_unsigned( 3850, 16)), --  3850 / 0x0f0a
    5414 => std_logic_vector(to_unsigned( 4422, 16)), --  4422 / 0x1146 -- last item of row
    5415 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5416 => std_logic_vector(to_unsigned( 5924, 16)), --  5924 / 0x1724
    5417 => std_logic_vector(to_unsigned(  290, 16)), --   290 / 0x0122 -- last item of row
    5418 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5419 => std_logic_vector(to_unsigned( 1467, 16)), --  1467 / 0x05bb
    5420 => std_logic_vector(to_unsigned( 4049, 16)), --  4049 / 0x0fd1 -- last item of row
    5421 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5422 => std_logic_vector(to_unsigned( 7820, 16)), --  7820 / 0x1e8c
    5423 => std_logic_vector(to_unsigned( 2242, 16)), --  2242 / 0x08c2 -- last item of row
    5424 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5425 => std_logic_vector(to_unsigned( 4606, 16)), --  4606 / 0x11fe
    5426 => std_logic_vector(to_unsigned( 3080, 16)), --  3080 / 0x0c08 -- last item of row
    5427 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5428 => std_logic_vector(to_unsigned( 4633, 16)), --  4633 / 0x1219
    5429 => std_logic_vector(to_unsigned( 7877, 16)), --  7877 / 0x1ec5 -- last item of row
    5430 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5431 => std_logic_vector(to_unsigned( 3884, 16)), --  3884 / 0x0f2c
    5432 => std_logic_vector(to_unsigned( 6868, 16)), --  6868 / 0x1ad4 -- last item of row
    5433 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5434 => std_logic_vector(to_unsigned( 8935, 16)), --  8935 / 0x22e7
    5435 => std_logic_vector(to_unsigned( 4996, 16)), --  4996 / 0x1384 -- last item of row
    5436 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5437 => std_logic_vector(to_unsigned( 3028, 16)), --  3028 / 0x0bd4
    5438 => std_logic_vector(to_unsigned(  764, 16)), --   764 / 0x02fc -- last item of row
    5439 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5440 => std_logic_vector(to_unsigned( 5988, 16)), --  5988 / 0x1764
    5441 => std_logic_vector(to_unsigned( 1057, 16)), --  1057 / 0x0421 -- last item of row
    5442 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5443 => std_logic_vector(to_unsigned( 7411, 16)), --  7411 / 0x1cf3
    5444 => std_logic_vector(to_unsigned( 3450, 16)), --  3450 / 0x0d7a -- last item of row
    -- Table for fecframe_short, C1_3
    5445 => std_logic_vector(to_unsigned(  416, 16)), --   416 / 0x01a0
    5446 => std_logic_vector(to_unsigned( 8909, 16)), --  8909 / 0x22cd
    5447 => std_logic_vector(to_unsigned( 4156, 16)), --  4156 / 0x103c
    5448 => std_logic_vector(to_unsigned( 3216, 16)), --  3216 / 0x0c90
    5449 => std_logic_vector(to_unsigned( 3112, 16)), --  3112 / 0x0c28
    5450 => std_logic_vector(to_unsigned( 2560, 16)), --  2560 / 0x0a00
    5451 => std_logic_vector(to_unsigned( 2912, 16)), --  2912 / 0x0b60
    5452 => std_logic_vector(to_unsigned( 6405, 16)), --  6405 / 0x1905
    5453 => std_logic_vector(to_unsigned( 8593, 16)), --  8593 / 0x2191
    5454 => std_logic_vector(to_unsigned( 4969, 16)), --  4969 / 0x1369
    5455 => std_logic_vector(to_unsigned( 6723, 16)), --  6723 / 0x1a43
    5456 => std_logic_vector(to_unsigned( 6912, 16)), --  6912 / 0x1b00 -- last item of row
    5457 => std_logic_vector(to_unsigned( 8978, 16)), --  8978 / 0x2312
    5458 => std_logic_vector(to_unsigned( 3011, 16)), --  3011 / 0x0bc3
    5459 => std_logic_vector(to_unsigned( 4339, 16)), --  4339 / 0x10f3
    5460 => std_logic_vector(to_unsigned( 9312, 16)), --  9312 / 0x2460
    5461 => std_logic_vector(to_unsigned( 6396, 16)), --  6396 / 0x18fc
    5462 => std_logic_vector(to_unsigned( 2957, 16)), --  2957 / 0x0b8d
    5463 => std_logic_vector(to_unsigned( 7288, 16)), --  7288 / 0x1c78
    5464 => std_logic_vector(to_unsigned( 5485, 16)), --  5485 / 0x156d
    5465 => std_logic_vector(to_unsigned( 6031, 16)), --  6031 / 0x178f
    5466 => std_logic_vector(to_unsigned(10218, 16)), -- 10218 / 0x27ea
    5467 => std_logic_vector(to_unsigned( 2226, 16)), --  2226 / 0x08b2
    5468 => std_logic_vector(to_unsigned( 3575, 16)), --  3575 / 0x0df7 -- last item of row
    5469 => std_logic_vector(to_unsigned( 3383, 16)), --  3383 / 0x0d37
    5470 => std_logic_vector(to_unsigned(10059, 16)), -- 10059 / 0x274b
    5471 => std_logic_vector(to_unsigned( 1114, 16)), --  1114 / 0x045a
    5472 => std_logic_vector(to_unsigned(10008, 16)), -- 10008 / 0x2718
    5473 => std_logic_vector(to_unsigned(10147, 16)), -- 10147 / 0x27a3
    5474 => std_logic_vector(to_unsigned( 9384, 16)), --  9384 / 0x24a8
    5475 => std_logic_vector(to_unsigned( 4290, 16)), --  4290 / 0x10c2
    5476 => std_logic_vector(to_unsigned(  434, 16)), --   434 / 0x01b2
    5477 => std_logic_vector(to_unsigned( 5139, 16)), --  5139 / 0x1413
    5478 => std_logic_vector(to_unsigned( 3536, 16)), --  3536 / 0x0dd0
    5479 => std_logic_vector(to_unsigned( 1965, 16)), --  1965 / 0x07ad
    5480 => std_logic_vector(to_unsigned( 2291, 16)), --  2291 / 0x08f3 -- last item of row
    5481 => std_logic_vector(to_unsigned( 2797, 16)), --  2797 / 0x0aed
    5482 => std_logic_vector(to_unsigned( 3693, 16)), --  3693 / 0x0e6d
    5483 => std_logic_vector(to_unsigned( 7615, 16)), --  7615 / 0x1dbf
    5484 => std_logic_vector(to_unsigned( 7077, 16)), --  7077 / 0x1ba5
    5485 => std_logic_vector(to_unsigned(  743, 16)), --   743 / 0x02e7
    5486 => std_logic_vector(to_unsigned( 1941, 16)), --  1941 / 0x0795
    5487 => std_logic_vector(to_unsigned( 8716, 16)), --  8716 / 0x220c
    5488 => std_logic_vector(to_unsigned( 6215, 16)), --  6215 / 0x1847
    5489 => std_logic_vector(to_unsigned( 3840, 16)), --  3840 / 0x0f00
    5490 => std_logic_vector(to_unsigned( 5140, 16)), --  5140 / 0x1414
    5491 => std_logic_vector(to_unsigned( 4582, 16)), --  4582 / 0x11e6
    5492 => std_logic_vector(to_unsigned( 5420, 16)), --  5420 / 0x152c -- last item of row
    5493 => std_logic_vector(to_unsigned( 6110, 16)), --  6110 / 0x17de
    5494 => std_logic_vector(to_unsigned( 8551, 16)), --  8551 / 0x2167
    5495 => std_logic_vector(to_unsigned( 1515, 16)), --  1515 / 0x05eb
    5496 => std_logic_vector(to_unsigned( 7404, 16)), --  7404 / 0x1cec
    5497 => std_logic_vector(to_unsigned( 4879, 16)), --  4879 / 0x130f
    5498 => std_logic_vector(to_unsigned( 4946, 16)), --  4946 / 0x1352
    5499 => std_logic_vector(to_unsigned( 5383, 16)), --  5383 / 0x1507
    5500 => std_logic_vector(to_unsigned( 1831, 16)), --  1831 / 0x0727
    5501 => std_logic_vector(to_unsigned( 3441, 16)), --  3441 / 0x0d71
    5502 => std_logic_vector(to_unsigned( 9569, 16)), --  9569 / 0x2561
    5503 => std_logic_vector(to_unsigned(10472, 16)), -- 10472 / 0x28e8
    5504 => std_logic_vector(to_unsigned( 4306, 16)), --  4306 / 0x10d2 -- last item of row
    5505 => std_logic_vector(to_unsigned( 1505, 16)), --  1505 / 0x05e1
    5506 => std_logic_vector(to_unsigned( 5682, 16)), --  5682 / 0x1632
    5507 => std_logic_vector(to_unsigned( 7778, 16)), --  7778 / 0x1e62 -- last item of row
    5508 => std_logic_vector(to_unsigned( 7172, 16)), --  7172 / 0x1c04
    5509 => std_logic_vector(to_unsigned( 6830, 16)), --  6830 / 0x1aae
    5510 => std_logic_vector(to_unsigned( 6623, 16)), --  6623 / 0x19df -- last item of row
    5511 => std_logic_vector(to_unsigned( 7281, 16)), --  7281 / 0x1c71
    5512 => std_logic_vector(to_unsigned( 3941, 16)), --  3941 / 0x0f65
    5513 => std_logic_vector(to_unsigned( 3505, 16)), --  3505 / 0x0db1 -- last item of row
    5514 => std_logic_vector(to_unsigned(10270, 16)), -- 10270 / 0x281e
    5515 => std_logic_vector(to_unsigned( 8669, 16)), --  8669 / 0x21dd
    5516 => std_logic_vector(to_unsigned(  914, 16)), --   914 / 0x0392 -- last item of row
    5517 => std_logic_vector(to_unsigned( 3622, 16)), --  3622 / 0x0e26
    5518 => std_logic_vector(to_unsigned( 7563, 16)), --  7563 / 0x1d8b
    5519 => std_logic_vector(to_unsigned( 9388, 16)), --  9388 / 0x24ac -- last item of row
    5520 => std_logic_vector(to_unsigned( 9930, 16)), --  9930 / 0x26ca
    5521 => std_logic_vector(to_unsigned( 5058, 16)), --  5058 / 0x13c2
    5522 => std_logic_vector(to_unsigned( 4554, 16)), --  4554 / 0x11ca -- last item of row
    5523 => std_logic_vector(to_unsigned( 4844, 16)), --  4844 / 0x12ec
    5524 => std_logic_vector(to_unsigned( 9609, 16)), --  9609 / 0x2589
    5525 => std_logic_vector(to_unsigned( 2707, 16)), --  2707 / 0x0a93 -- last item of row
    5526 => std_logic_vector(to_unsigned( 6883, 16)), --  6883 / 0x1ae3
    5527 => std_logic_vector(to_unsigned( 3237, 16)), --  3237 / 0x0ca5
    5528 => std_logic_vector(to_unsigned( 1714, 16)), --  1714 / 0x06b2 -- last item of row
    5529 => std_logic_vector(to_unsigned( 4768, 16)), --  4768 / 0x12a0
    5530 => std_logic_vector(to_unsigned( 3878, 16)), --  3878 / 0x0f26
    5531 => std_logic_vector(to_unsigned(10017, 16)), -- 10017 / 0x2721 -- last item of row
    5532 => std_logic_vector(to_unsigned(10127, 16)), -- 10127 / 0x278f
    5533 => std_logic_vector(to_unsigned( 3334, 16)), --  3334 / 0x0d06
    5534 => std_logic_vector(to_unsigned( 8267, 16)), --  8267 / 0x204b -- last item of row
    -- Table for fecframe_short, C1_4
    5535 => std_logic_vector(to_unsigned( 6295, 16)), --  6295 / 0x1897
    5536 => std_logic_vector(to_unsigned( 9626, 16)), --  9626 / 0x259a
    5537 => std_logic_vector(to_unsigned(  304, 16)), --   304 / 0x0130
    5538 => std_logic_vector(to_unsigned( 7695, 16)), --  7695 / 0x1e0f
    5539 => std_logic_vector(to_unsigned( 4839, 16)), --  4839 / 0x12e7
    5540 => std_logic_vector(to_unsigned( 4936, 16)), --  4936 / 0x1348
    5541 => std_logic_vector(to_unsigned( 1660, 16)), --  1660 / 0x067c
    5542 => std_logic_vector(to_unsigned(  144, 16)), --   144 / 0x0090
    5543 => std_logic_vector(to_unsigned(11203, 16)), -- 11203 / 0x2bc3
    5544 => std_logic_vector(to_unsigned( 5567, 16)), --  5567 / 0x15bf
    5545 => std_logic_vector(to_unsigned( 6347, 16)), --  6347 / 0x18cb
    5546 => std_logic_vector(to_unsigned(12557, 16)), -- 12557 / 0x310d -- last item of row
    5547 => std_logic_vector(to_unsigned(10691, 16)), -- 10691 / 0x29c3
    5548 => std_logic_vector(to_unsigned( 4988, 16)), --  4988 / 0x137c
    5549 => std_logic_vector(to_unsigned( 3859, 16)), --  3859 / 0x0f13
    5550 => std_logic_vector(to_unsigned( 3734, 16)), --  3734 / 0x0e96
    5551 => std_logic_vector(to_unsigned( 3071, 16)), --  3071 / 0x0bff
    5552 => std_logic_vector(to_unsigned( 3494, 16)), --  3494 / 0x0da6
    5553 => std_logic_vector(to_unsigned( 7687, 16)), --  7687 / 0x1e07
    5554 => std_logic_vector(to_unsigned(10313, 16)), -- 10313 / 0x2849
    5555 => std_logic_vector(to_unsigned( 5964, 16)), --  5964 / 0x174c
    5556 => std_logic_vector(to_unsigned( 8069, 16)), --  8069 / 0x1f85
    5557 => std_logic_vector(to_unsigned( 8296, 16)), --  8296 / 0x2068
    5558 => std_logic_vector(to_unsigned(11090, 16)), -- 11090 / 0x2b52 -- last item of row
    5559 => std_logic_vector(to_unsigned(10774, 16)), -- 10774 / 0x2a16
    5560 => std_logic_vector(to_unsigned( 3613, 16)), --  3613 / 0x0e1d
    5561 => std_logic_vector(to_unsigned( 5208, 16)), --  5208 / 0x1458
    5562 => std_logic_vector(to_unsigned(11177, 16)), -- 11177 / 0x2ba9
    5563 => std_logic_vector(to_unsigned( 7676, 16)), --  7676 / 0x1dfc
    5564 => std_logic_vector(to_unsigned( 3549, 16)), --  3549 / 0x0ddd
    5565 => std_logic_vector(to_unsigned( 8746, 16)), --  8746 / 0x222a
    5566 => std_logic_vector(to_unsigned( 6583, 16)), --  6583 / 0x19b7
    5567 => std_logic_vector(to_unsigned( 7239, 16)), --  7239 / 0x1c47
    5568 => std_logic_vector(to_unsigned(12265, 16)), -- 12265 / 0x2fe9
    5569 => std_logic_vector(to_unsigned( 2674, 16)), --  2674 / 0x0a72
    5570 => std_logic_vector(to_unsigned( 4292, 16)), --  4292 / 0x10c4 -- last item of row
    5571 => std_logic_vector(to_unsigned(11869, 16)), -- 11869 / 0x2e5d
    5572 => std_logic_vector(to_unsigned( 3708, 16)), --  3708 / 0x0e7c
    5573 => std_logic_vector(to_unsigned( 5981, 16)), --  5981 / 0x175d
    5574 => std_logic_vector(to_unsigned( 8718, 16)), --  8718 / 0x220e
    5575 => std_logic_vector(to_unsigned( 4908, 16)), --  4908 / 0x132c
    5576 => std_logic_vector(to_unsigned(10650, 16)), -- 10650 / 0x299a
    5577 => std_logic_vector(to_unsigned( 6805, 16)), --  6805 / 0x1a95
    5578 => std_logic_vector(to_unsigned( 3334, 16)), --  3334 / 0x0d06
    5579 => std_logic_vector(to_unsigned( 2627, 16)), --  2627 / 0x0a43
    5580 => std_logic_vector(to_unsigned(10461, 16)), -- 10461 / 0x28dd
    5581 => std_logic_vector(to_unsigned( 9285, 16)), --  9285 / 0x2445
    5582 => std_logic_vector(to_unsigned(11120, 16)), -- 11120 / 0x2b70 -- last item of row
    5583 => std_logic_vector(to_unsigned( 7844, 16)), --  7844 / 0x1ea4
    5584 => std_logic_vector(to_unsigned( 3079, 16)), --  3079 / 0x0c07
    5585 => std_logic_vector(to_unsigned(10773, 16)), -- 10773 / 0x2a15 -- last item of row
    5586 => std_logic_vector(to_unsigned( 3385, 16)), --  3385 / 0x0d39
    5587 => std_logic_vector(to_unsigned(10854, 16)), -- 10854 / 0x2a66
    5588 => std_logic_vector(to_unsigned( 5747, 16)), --  5747 / 0x1673 -- last item of row
    5589 => std_logic_vector(to_unsigned( 1360, 16)), --  1360 / 0x0550
    5590 => std_logic_vector(to_unsigned(12010, 16)), -- 12010 / 0x2eea
    5591 => std_logic_vector(to_unsigned(12202, 16)), -- 12202 / 0x2faa -- last item of row
    5592 => std_logic_vector(to_unsigned( 6189, 16)), --  6189 / 0x182d
    5593 => std_logic_vector(to_unsigned( 4241, 16)), --  4241 / 0x1091
    5594 => std_logic_vector(to_unsigned( 2343, 16)), --  2343 / 0x0927 -- last item of row
    5595 => std_logic_vector(to_unsigned( 9840, 16)), --  9840 / 0x2670
    5596 => std_logic_vector(to_unsigned(12726, 16)), -- 12726 / 0x31b6
    5597 => std_logic_vector(to_unsigned( 4977, 16)), --  4977 / 0x1371 -- last item of row
    -- Table for fecframe_short, C2_3
    5598 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5599 => std_logic_vector(to_unsigned( 2084, 16)), --  2084 / 0x0824
    5600 => std_logic_vector(to_unsigned( 1613, 16)), --  1613 / 0x064d
    5601 => std_logic_vector(to_unsigned( 1548, 16)), --  1548 / 0x060c
    5602 => std_logic_vector(to_unsigned( 1286, 16)), --  1286 / 0x0506
    5603 => std_logic_vector(to_unsigned( 1460, 16)), --  1460 / 0x05b4
    5604 => std_logic_vector(to_unsigned( 3196, 16)), --  3196 / 0x0c7c
    5605 => std_logic_vector(to_unsigned( 4297, 16)), --  4297 / 0x10c9
    5606 => std_logic_vector(to_unsigned( 2481, 16)), --  2481 / 0x09b1
    5607 => std_logic_vector(to_unsigned( 3369, 16)), --  3369 / 0x0d29
    5608 => std_logic_vector(to_unsigned( 3451, 16)), --  3451 / 0x0d7b
    5609 => std_logic_vector(to_unsigned( 4620, 16)), --  4620 / 0x120c
    5610 => std_logic_vector(to_unsigned( 2622, 16)), --  2622 / 0x0a3e -- last item of row
    5611 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5612 => std_logic_vector(to_unsigned(  122, 16)), --   122 / 0x007a
    5613 => std_logic_vector(to_unsigned( 1516, 16)), --  1516 / 0x05ec
    5614 => std_logic_vector(to_unsigned( 3448, 16)), --  3448 / 0x0d78
    5615 => std_logic_vector(to_unsigned( 2880, 16)), --  2880 / 0x0b40
    5616 => std_logic_vector(to_unsigned( 1407, 16)), --  1407 / 0x057f
    5617 => std_logic_vector(to_unsigned( 1847, 16)), --  1847 / 0x0737
    5618 => std_logic_vector(to_unsigned( 3799, 16)), --  3799 / 0x0ed7
    5619 => std_logic_vector(to_unsigned( 3529, 16)), --  3529 / 0x0dc9
    5620 => std_logic_vector(to_unsigned(  373, 16)), --   373 / 0x0175
    5621 => std_logic_vector(to_unsigned(  971, 16)), --   971 / 0x03cb
    5622 => std_logic_vector(to_unsigned( 4358, 16)), --  4358 / 0x1106
    5623 => std_logic_vector(to_unsigned( 3108, 16)), --  3108 / 0x0c24 -- last item of row
    5624 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5625 => std_logic_vector(to_unsigned(  259, 16)), --   259 / 0x0103
    5626 => std_logic_vector(to_unsigned( 3399, 16)), --  3399 / 0x0d47
    5627 => std_logic_vector(to_unsigned(  929, 16)), --   929 / 0x03a1
    5628 => std_logic_vector(to_unsigned( 2650, 16)), --  2650 / 0x0a5a
    5629 => std_logic_vector(to_unsigned(  864, 16)), --   864 / 0x0360
    5630 => std_logic_vector(to_unsigned( 3996, 16)), --  3996 / 0x0f9c
    5631 => std_logic_vector(to_unsigned( 3833, 16)), --  3833 / 0x0ef9
    5632 => std_logic_vector(to_unsigned(  107, 16)), --   107 / 0x006b
    5633 => std_logic_vector(to_unsigned( 5287, 16)), --  5287 / 0x14a7
    5634 => std_logic_vector(to_unsigned(  164, 16)), --   164 / 0x00a4
    5635 => std_logic_vector(to_unsigned( 3125, 16)), --  3125 / 0x0c35
    5636 => std_logic_vector(to_unsigned( 2350, 16)), --  2350 / 0x092e -- last item of row
    5637 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5638 => std_logic_vector(to_unsigned(  342, 16)), --   342 / 0x0156
    5639 => std_logic_vector(to_unsigned( 3529, 16)), --  3529 / 0x0dc9 -- last item of row
    5640 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5641 => std_logic_vector(to_unsigned( 4198, 16)), --  4198 / 0x1066
    5642 => std_logic_vector(to_unsigned( 2147, 16)), --  2147 / 0x0863 -- last item of row
    5643 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5644 => std_logic_vector(to_unsigned( 1880, 16)), --  1880 / 0x0758
    5645 => std_logic_vector(to_unsigned( 4836, 16)), --  4836 / 0x12e4 -- last item of row
    5646 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5647 => std_logic_vector(to_unsigned( 3864, 16)), --  3864 / 0x0f18
    5648 => std_logic_vector(to_unsigned( 4910, 16)), --  4910 / 0x132e -- last item of row
    5649 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5650 => std_logic_vector(to_unsigned(  243, 16)), --   243 / 0x00f3
    5651 => std_logic_vector(to_unsigned( 1542, 16)), --  1542 / 0x0606 -- last item of row
    5652 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5653 => std_logic_vector(to_unsigned( 3011, 16)), --  3011 / 0x0bc3
    5654 => std_logic_vector(to_unsigned( 1436, 16)), --  1436 / 0x059c -- last item of row
    5655 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5656 => std_logic_vector(to_unsigned( 2167, 16)), --  2167 / 0x0877
    5657 => std_logic_vector(to_unsigned( 2512, 16)), --  2512 / 0x09d0 -- last item of row
    5658 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5659 => std_logic_vector(to_unsigned( 4606, 16)), --  4606 / 0x11fe
    5660 => std_logic_vector(to_unsigned( 1003, 16)), --  1003 / 0x03eb -- last item of row
    5661 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5662 => std_logic_vector(to_unsigned( 2835, 16)), --  2835 / 0x0b13
    5663 => std_logic_vector(to_unsigned(  705, 16)), --   705 / 0x02c1 -- last item of row
    5664 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5665 => std_logic_vector(to_unsigned( 3426, 16)), --  3426 / 0x0d62
    5666 => std_logic_vector(to_unsigned( 2365, 16)), --  2365 / 0x093d -- last item of row
    5667 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5668 => std_logic_vector(to_unsigned( 3848, 16)), --  3848 / 0x0f08
    5669 => std_logic_vector(to_unsigned( 2474, 16)), --  2474 / 0x09aa -- last item of row
    5670 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5671 => std_logic_vector(to_unsigned( 1360, 16)), --  1360 / 0x0550
    5672 => std_logic_vector(to_unsigned( 1743, 16)), --  1743 / 0x06cf -- last item of row
    5673 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5674 => std_logic_vector(to_unsigned(  163, 16)), --   163 / 0x00a3
    5675 => std_logic_vector(to_unsigned( 2536, 16)), --  2536 / 0x09e8 -- last item of row
    5676 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5677 => std_logic_vector(to_unsigned( 2583, 16)), --  2583 / 0x0a17
    5678 => std_logic_vector(to_unsigned( 1180, 16)), --  1180 / 0x049c -- last item of row
    5679 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5680 => std_logic_vector(to_unsigned( 1542, 16)), --  1542 / 0x0606
    5681 => std_logic_vector(to_unsigned(  509, 16)), --   509 / 0x01fd -- last item of row
    5682 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5683 => std_logic_vector(to_unsigned( 4418, 16)), --  4418 / 0x1142
    5684 => std_logic_vector(to_unsigned( 1005, 16)), --  1005 / 0x03ed -- last item of row
    5685 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5686 => std_logic_vector(to_unsigned( 5212, 16)), --  5212 / 0x145c
    5687 => std_logic_vector(to_unsigned( 5117, 16)), --  5117 / 0x13fd -- last item of row
    5688 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5689 => std_logic_vector(to_unsigned( 2155, 16)), --  2155 / 0x086b
    5690 => std_logic_vector(to_unsigned( 2922, 16)), --  2922 / 0x0b6a -- last item of row
    5691 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5692 => std_logic_vector(to_unsigned(  347, 16)), --   347 / 0x015b
    5693 => std_logic_vector(to_unsigned( 2696, 16)), --  2696 / 0x0a88 -- last item of row
    5694 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5695 => std_logic_vector(to_unsigned(  226, 16)), --   226 / 0x00e2
    5696 => std_logic_vector(to_unsigned( 4296, 16)), --  4296 / 0x10c8 -- last item of row
    5697 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5698 => std_logic_vector(to_unsigned( 1560, 16)), --  1560 / 0x0618
    5699 => std_logic_vector(to_unsigned(  487, 16)), --   487 / 0x01e7 -- last item of row
    5700 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5701 => std_logic_vector(to_unsigned( 3926, 16)), --  3926 / 0x0f56
    5702 => std_logic_vector(to_unsigned( 1640, 16)), --  1640 / 0x0668 -- last item of row
    5703 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5704 => std_logic_vector(to_unsigned(  149, 16)), --   149 / 0x0095
    5705 => std_logic_vector(to_unsigned( 2928, 16)), --  2928 / 0x0b70 -- last item of row
    5706 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5707 => std_logic_vector(to_unsigned( 2364, 16)), --  2364 / 0x093c
    5708 => std_logic_vector(to_unsigned(  563, 16)), --   563 / 0x0233 -- last item of row
    5709 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    5710 => std_logic_vector(to_unsigned(  635, 16)), --   635 / 0x027b
    5711 => std_logic_vector(to_unsigned(  688, 16)), --   688 / 0x02b0 -- last item of row
    5712 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    5713 => std_logic_vector(to_unsigned(  231, 16)), --   231 / 0x00e7
    5714 => std_logic_vector(to_unsigned( 1684, 16)), --  1684 / 0x0694 -- last item of row
    5715 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    5716 => std_logic_vector(to_unsigned( 1129, 16)), --  1129 / 0x0469
    5717 => std_logic_vector(to_unsigned( 3894, 16)), --  3894 / 0x0f36 -- last item of row
    -- Table for fecframe_short, C2_5
    5718 => std_logic_vector(to_unsigned( 5650, 16)), --  5650 / 0x1612
    5719 => std_logic_vector(to_unsigned( 4143, 16)), --  4143 / 0x102f
    5720 => std_logic_vector(to_unsigned( 8750, 16)), --  8750 / 0x222e
    5721 => std_logic_vector(to_unsigned(  583, 16)), --   583 / 0x0247
    5722 => std_logic_vector(to_unsigned( 6720, 16)), --  6720 / 0x1a40
    5723 => std_logic_vector(to_unsigned( 8071, 16)), --  8071 / 0x1f87
    5724 => std_logic_vector(to_unsigned(  635, 16)), --   635 / 0x027b
    5725 => std_logic_vector(to_unsigned( 1767, 16)), --  1767 / 0x06e7
    5726 => std_logic_vector(to_unsigned( 1344, 16)), --  1344 / 0x0540
    5727 => std_logic_vector(to_unsigned( 6922, 16)), --  6922 / 0x1b0a
    5728 => std_logic_vector(to_unsigned(  738, 16)), --   738 / 0x02e2
    5729 => std_logic_vector(to_unsigned( 6658, 16)), --  6658 / 0x1a02 -- last item of row
    5730 => std_logic_vector(to_unsigned( 5696, 16)), --  5696 / 0x1640
    5731 => std_logic_vector(to_unsigned( 1685, 16)), --  1685 / 0x0695
    5732 => std_logic_vector(to_unsigned( 3207, 16)), --  3207 / 0x0c87
    5733 => std_logic_vector(to_unsigned(  415, 16)), --   415 / 0x019f
    5734 => std_logic_vector(to_unsigned( 7019, 16)), --  7019 / 0x1b6b
    5735 => std_logic_vector(to_unsigned( 5023, 16)), --  5023 / 0x139f
    5736 => std_logic_vector(to_unsigned( 5608, 16)), --  5608 / 0x15e8
    5737 => std_logic_vector(to_unsigned( 2605, 16)), --  2605 / 0x0a2d
    5738 => std_logic_vector(to_unsigned(  857, 16)), --   857 / 0x0359
    5739 => std_logic_vector(to_unsigned( 6915, 16)), --  6915 / 0x1b03
    5740 => std_logic_vector(to_unsigned( 1770, 16)), --  1770 / 0x06ea
    5741 => std_logic_vector(to_unsigned( 8016, 16)), --  8016 / 0x1f50 -- last item of row
    5742 => std_logic_vector(to_unsigned( 3992, 16)), --  3992 / 0x0f98
    5743 => std_logic_vector(to_unsigned(  771, 16)), --   771 / 0x0303
    5744 => std_logic_vector(to_unsigned( 2190, 16)), --  2190 / 0x088e
    5745 => std_logic_vector(to_unsigned( 7258, 16)), --  7258 / 0x1c5a
    5746 => std_logic_vector(to_unsigned( 8970, 16)), --  8970 / 0x230a
    5747 => std_logic_vector(to_unsigned( 7792, 16)), --  7792 / 0x1e70
    5748 => std_logic_vector(to_unsigned( 1802, 16)), --  1802 / 0x070a
    5749 => std_logic_vector(to_unsigned( 1866, 16)), --  1866 / 0x074a
    5750 => std_logic_vector(to_unsigned( 6137, 16)), --  6137 / 0x17f9
    5751 => std_logic_vector(to_unsigned( 8841, 16)), --  8841 / 0x2289
    5752 => std_logic_vector(to_unsigned(  886, 16)), --   886 / 0x0376
    5753 => std_logic_vector(to_unsigned( 1931, 16)), --  1931 / 0x078b -- last item of row
    5754 => std_logic_vector(to_unsigned( 4108, 16)), --  4108 / 0x100c
    5755 => std_logic_vector(to_unsigned( 3781, 16)), --  3781 / 0x0ec5
    5756 => std_logic_vector(to_unsigned( 7577, 16)), --  7577 / 0x1d99
    5757 => std_logic_vector(to_unsigned( 6810, 16)), --  6810 / 0x1a9a
    5758 => std_logic_vector(to_unsigned( 9322, 16)), --  9322 / 0x246a
    5759 => std_logic_vector(to_unsigned( 8226, 16)), --  8226 / 0x2022
    5760 => std_logic_vector(to_unsigned( 5396, 16)), --  5396 / 0x1514
    5761 => std_logic_vector(to_unsigned( 5867, 16)), --  5867 / 0x16eb
    5762 => std_logic_vector(to_unsigned( 4428, 16)), --  4428 / 0x114c
    5763 => std_logic_vector(to_unsigned( 8827, 16)), --  8827 / 0x227b
    5764 => std_logic_vector(to_unsigned( 7766, 16)), --  7766 / 0x1e56
    5765 => std_logic_vector(to_unsigned( 2254, 16)), --  2254 / 0x08ce -- last item of row
    5766 => std_logic_vector(to_unsigned( 4247, 16)), --  4247 / 0x1097
    5767 => std_logic_vector(to_unsigned(  888, 16)), --   888 / 0x0378
    5768 => std_logic_vector(to_unsigned( 4367, 16)), --  4367 / 0x110f
    5769 => std_logic_vector(to_unsigned( 8821, 16)), --  8821 / 0x2275
    5770 => std_logic_vector(to_unsigned( 9660, 16)), --  9660 / 0x25bc
    5771 => std_logic_vector(to_unsigned(  324, 16)), --   324 / 0x0144
    5772 => std_logic_vector(to_unsigned( 5864, 16)), --  5864 / 0x16e8
    5773 => std_logic_vector(to_unsigned( 4774, 16)), --  4774 / 0x12a6
    5774 => std_logic_vector(to_unsigned(  227, 16)), --   227 / 0x00e3
    5775 => std_logic_vector(to_unsigned( 7889, 16)), --  7889 / 0x1ed1
    5776 => std_logic_vector(to_unsigned( 6405, 16)), --  6405 / 0x1905
    5777 => std_logic_vector(to_unsigned( 8963, 16)), --  8963 / 0x2303 -- last item of row
    5778 => std_logic_vector(to_unsigned( 9693, 16)), --  9693 / 0x25dd
    5779 => std_logic_vector(to_unsigned(  500, 16)), --   500 / 0x01f4
    5780 => std_logic_vector(to_unsigned( 2520, 16)), --  2520 / 0x09d8
    5781 => std_logic_vector(to_unsigned( 2227, 16)), --  2227 / 0x08b3
    5782 => std_logic_vector(to_unsigned( 1811, 16)), --  1811 / 0x0713
    5783 => std_logic_vector(to_unsigned( 9330, 16)), --  9330 / 0x2472
    5784 => std_logic_vector(to_unsigned( 1928, 16)), --  1928 / 0x0788
    5785 => std_logic_vector(to_unsigned( 5140, 16)), --  5140 / 0x1414
    5786 => std_logic_vector(to_unsigned( 4030, 16)), --  4030 / 0x0fbe
    5787 => std_logic_vector(to_unsigned( 4824, 16)), --  4824 / 0x12d8
    5788 => std_logic_vector(to_unsigned(  806, 16)), --   806 / 0x0326
    5789 => std_logic_vector(to_unsigned( 3134, 16)), --  3134 / 0x0c3e -- last item of row
    5790 => std_logic_vector(to_unsigned( 1652, 16)), --  1652 / 0x0674
    5791 => std_logic_vector(to_unsigned( 8171, 16)), --  8171 / 0x1feb
    5792 => std_logic_vector(to_unsigned( 1435, 16)), --  1435 / 0x059b -- last item of row
    5793 => std_logic_vector(to_unsigned( 3366, 16)), --  3366 / 0x0d26
    5794 => std_logic_vector(to_unsigned( 6543, 16)), --  6543 / 0x198f
    5795 => std_logic_vector(to_unsigned( 3745, 16)), --  3745 / 0x0ea1 -- last item of row
    5796 => std_logic_vector(to_unsigned( 9286, 16)), --  9286 / 0x2446
    5797 => std_logic_vector(to_unsigned( 8509, 16)), --  8509 / 0x213d
    5798 => std_logic_vector(to_unsigned( 4645, 16)), --  4645 / 0x1225 -- last item of row
    5799 => std_logic_vector(to_unsigned( 7397, 16)), --  7397 / 0x1ce5
    5800 => std_logic_vector(to_unsigned( 5790, 16)), --  5790 / 0x169e
    5801 => std_logic_vector(to_unsigned( 8972, 16)), --  8972 / 0x230c -- last item of row
    5802 => std_logic_vector(to_unsigned( 6597, 16)), --  6597 / 0x19c5
    5803 => std_logic_vector(to_unsigned( 4422, 16)), --  4422 / 0x1146
    5804 => std_logic_vector(to_unsigned( 1799, 16)), --  1799 / 0x0707 -- last item of row
    5805 => std_logic_vector(to_unsigned( 9276, 16)), --  9276 / 0x243c
    5806 => std_logic_vector(to_unsigned( 4041, 16)), --  4041 / 0x0fc9
    5807 => std_logic_vector(to_unsigned( 3847, 16)), --  3847 / 0x0f07 -- last item of row
    5808 => std_logic_vector(to_unsigned( 8683, 16)), --  8683 / 0x21eb
    5809 => std_logic_vector(to_unsigned( 7378, 16)), --  7378 / 0x1cd2
    5810 => std_logic_vector(to_unsigned( 4946, 16)), --  4946 / 0x1352 -- last item of row
    5811 => std_logic_vector(to_unsigned( 5348, 16)), --  5348 / 0x14e4
    5812 => std_logic_vector(to_unsigned( 1993, 16)), --  1993 / 0x07c9
    5813 => std_logic_vector(to_unsigned( 9186, 16)), --  9186 / 0x23e2 -- last item of row
    5814 => std_logic_vector(to_unsigned( 6724, 16)), --  6724 / 0x1a44
    5815 => std_logic_vector(to_unsigned( 9015, 16)), --  9015 / 0x2337
    5816 => std_logic_vector(to_unsigned( 5646, 16)), --  5646 / 0x160e -- last item of row
    5817 => std_logic_vector(to_unsigned( 4502, 16)), --  4502 / 0x1196
    5818 => std_logic_vector(to_unsigned( 4439, 16)), --  4439 / 0x1157
    5819 => std_logic_vector(to_unsigned( 8474, 16)), --  8474 / 0x211a -- last item of row
    5820 => std_logic_vector(to_unsigned( 5107, 16)), --  5107 / 0x13f3
    5821 => std_logic_vector(to_unsigned( 7342, 16)), --  7342 / 0x1cae
    5822 => std_logic_vector(to_unsigned( 9442, 16)), --  9442 / 0x24e2 -- last item of row
    5823 => std_logic_vector(to_unsigned( 1387, 16)), --  1387 / 0x056b
    5824 => std_logic_vector(to_unsigned( 8910, 16)), --  8910 / 0x22ce
    5825 => std_logic_vector(to_unsigned( 2660, 16)), --  2660 / 0x0a64 -- last item of row
    -- Table for fecframe_short, C3_4
    5826 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5827 => std_logic_vector(to_unsigned( 3198, 16)), --  3198 / 0x0c7e
    5828 => std_logic_vector(to_unsigned(  478, 16)), --   478 / 0x01de
    5829 => std_logic_vector(to_unsigned( 4207, 16)), --  4207 / 0x106f
    5830 => std_logic_vector(to_unsigned( 1481, 16)), --  1481 / 0x05c9
    5831 => std_logic_vector(to_unsigned( 1009, 16)), --  1009 / 0x03f1
    5832 => std_logic_vector(to_unsigned( 2616, 16)), --  2616 / 0x0a38
    5833 => std_logic_vector(to_unsigned( 1924, 16)), --  1924 / 0x0784
    5834 => std_logic_vector(to_unsigned( 3437, 16)), --  3437 / 0x0d6d
    5835 => std_logic_vector(to_unsigned(  554, 16)), --   554 / 0x022a
    5836 => std_logic_vector(to_unsigned(  683, 16)), --   683 / 0x02ab
    5837 => std_logic_vector(to_unsigned( 1801, 16)), --  1801 / 0x0709 -- last item of row
    5838 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5839 => std_logic_vector(to_unsigned( 2681, 16)), --  2681 / 0x0a79
    5840 => std_logic_vector(to_unsigned( 2135, 16)), --  2135 / 0x0857 -- last item of row
    5841 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5842 => std_logic_vector(to_unsigned( 3107, 16)), --  3107 / 0x0c23
    5843 => std_logic_vector(to_unsigned( 4027, 16)), --  4027 / 0x0fbb -- last item of row
    5844 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5845 => std_logic_vector(to_unsigned( 2637, 16)), --  2637 / 0x0a4d
    5846 => std_logic_vector(to_unsigned( 3373, 16)), --  3373 / 0x0d2d -- last item of row
    5847 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5848 => std_logic_vector(to_unsigned( 3830, 16)), --  3830 / 0x0ef6
    5849 => std_logic_vector(to_unsigned( 3449, 16)), --  3449 / 0x0d79 -- last item of row
    5850 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5851 => std_logic_vector(to_unsigned( 4129, 16)), --  4129 / 0x1021
    5852 => std_logic_vector(to_unsigned( 2060, 16)), --  2060 / 0x080c -- last item of row
    5853 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5854 => std_logic_vector(to_unsigned( 4184, 16)), --  4184 / 0x1058
    5855 => std_logic_vector(to_unsigned( 2742, 16)), --  2742 / 0x0ab6 -- last item of row
    5856 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5857 => std_logic_vector(to_unsigned( 3946, 16)), --  3946 / 0x0f6a
    5858 => std_logic_vector(to_unsigned( 1070, 16)), --  1070 / 0x042e -- last item of row
    5859 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5860 => std_logic_vector(to_unsigned( 2239, 16)), --  2239 / 0x08bf
    5861 => std_logic_vector(to_unsigned(  984, 16)), --   984 / 0x03d8 -- last item of row
    5862 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5863 => std_logic_vector(to_unsigned( 1458, 16)), --  1458 / 0x05b2
    5864 => std_logic_vector(to_unsigned( 3031, 16)), --  3031 / 0x0bd7 -- last item of row
    5865 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5866 => std_logic_vector(to_unsigned( 3003, 16)), --  3003 / 0x0bbb
    5867 => std_logic_vector(to_unsigned( 1328, 16)), --  1328 / 0x0530 -- last item of row
    5868 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5869 => std_logic_vector(to_unsigned( 1137, 16)), --  1137 / 0x0471
    5870 => std_logic_vector(to_unsigned( 1716, 16)), --  1716 / 0x06b4 -- last item of row
    5871 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5872 => std_logic_vector(to_unsigned(  132, 16)), --   132 / 0x0084
    5873 => std_logic_vector(to_unsigned( 3725, 16)), --  3725 / 0x0e8d -- last item of row
    5874 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5875 => std_logic_vector(to_unsigned( 1817, 16)), --  1817 / 0x0719
    5876 => std_logic_vector(to_unsigned(  638, 16)), --   638 / 0x027e -- last item of row
    5877 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5878 => std_logic_vector(to_unsigned( 1774, 16)), --  1774 / 0x06ee
    5879 => std_logic_vector(to_unsigned( 3447, 16)), --  3447 / 0x0d77 -- last item of row
    5880 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5881 => std_logic_vector(to_unsigned( 3632, 16)), --  3632 / 0x0e30
    5882 => std_logic_vector(to_unsigned( 1257, 16)), --  1257 / 0x04e9 -- last item of row
    5883 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5884 => std_logic_vector(to_unsigned(  542, 16)), --   542 / 0x021e
    5885 => std_logic_vector(to_unsigned( 3694, 16)), --  3694 / 0x0e6e -- last item of row
    5886 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5887 => std_logic_vector(to_unsigned( 1015, 16)), --  1015 / 0x03f7
    5888 => std_logic_vector(to_unsigned( 1945, 16)), --  1945 / 0x0799 -- last item of row
    5889 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5890 => std_logic_vector(to_unsigned( 1948, 16)), --  1948 / 0x079c
    5891 => std_logic_vector(to_unsigned(  412, 16)), --   412 / 0x019c -- last item of row
    5892 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5893 => std_logic_vector(to_unsigned(  995, 16)), --   995 / 0x03e3
    5894 => std_logic_vector(to_unsigned( 2238, 16)), --  2238 / 0x08be -- last item of row
    5895 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5896 => std_logic_vector(to_unsigned( 4141, 16)), --  4141 / 0x102d
    5897 => std_logic_vector(to_unsigned( 1907, 16)), --  1907 / 0x0773 -- last item of row
    5898 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    5899 => std_logic_vector(to_unsigned( 2480, 16)), --  2480 / 0x09b0
    5900 => std_logic_vector(to_unsigned( 3079, 16)), --  3079 / 0x0c07 -- last item of row
    5901 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    5902 => std_logic_vector(to_unsigned( 3021, 16)), --  3021 / 0x0bcd
    5903 => std_logic_vector(to_unsigned( 1088, 16)), --  1088 / 0x0440 -- last item of row
    5904 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    5905 => std_logic_vector(to_unsigned(  713, 16)), --   713 / 0x02c9
    5906 => std_logic_vector(to_unsigned( 1379, 16)), --  1379 / 0x0563 -- last item of row
    5907 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    5908 => std_logic_vector(to_unsigned(  997, 16)), --   997 / 0x03e5
    5909 => std_logic_vector(to_unsigned( 3903, 16)), --  3903 / 0x0f3f -- last item of row
    5910 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    5911 => std_logic_vector(to_unsigned( 2323, 16)), --  2323 / 0x0913
    5912 => std_logic_vector(to_unsigned( 3361, 16)), --  3361 / 0x0d21 -- last item of row
    5913 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    5914 => std_logic_vector(to_unsigned( 1110, 16)), --  1110 / 0x0456
    5915 => std_logic_vector(to_unsigned(  986, 16)), --   986 / 0x03da -- last item of row
    5916 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    5917 => std_logic_vector(to_unsigned( 2532, 16)), --  2532 / 0x09e4
    5918 => std_logic_vector(to_unsigned(  142, 16)), --   142 / 0x008e -- last item of row
    5919 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    5920 => std_logic_vector(to_unsigned( 1690, 16)), --  1690 / 0x069a
    5921 => std_logic_vector(to_unsigned( 2405, 16)), --  2405 / 0x0965 -- last item of row
    5922 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    5923 => std_logic_vector(to_unsigned( 1298, 16)), --  1298 / 0x0512
    5924 => std_logic_vector(to_unsigned( 1881, 16)), --  1881 / 0x0759 -- last item of row
    5925 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    5926 => std_logic_vector(to_unsigned(  615, 16)), --   615 / 0x0267
    5927 => std_logic_vector(to_unsigned(  174, 16)), --   174 / 0x00ae -- last item of row
    5928 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    5929 => std_logic_vector(to_unsigned( 1648, 16)), --  1648 / 0x0670
    5930 => std_logic_vector(to_unsigned( 3112, 16)), --  3112 / 0x0c28 -- last item of row
    5931 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    5932 => std_logic_vector(to_unsigned( 1415, 16)), --  1415 / 0x0587
    5933 => std_logic_vector(to_unsigned( 2808, 16)), --  2808 / 0x0af8 -- last item of row
    -- Table for fecframe_short, C3_5
    5934 => std_logic_vector(to_unsigned( 2765, 16)), --  2765 / 0x0acd
    5935 => std_logic_vector(to_unsigned( 5713, 16)), --  5713 / 0x1651
    5936 => std_logic_vector(to_unsigned( 6426, 16)), --  6426 / 0x191a
    5937 => std_logic_vector(to_unsigned( 3596, 16)), --  3596 / 0x0e0c
    5938 => std_logic_vector(to_unsigned( 1374, 16)), --  1374 / 0x055e
    5939 => std_logic_vector(to_unsigned( 4811, 16)), --  4811 / 0x12cb
    5940 => std_logic_vector(to_unsigned( 2182, 16)), --  2182 / 0x0886
    5941 => std_logic_vector(to_unsigned(  544, 16)), --   544 / 0x0220
    5942 => std_logic_vector(to_unsigned( 3394, 16)), --  3394 / 0x0d42
    5943 => std_logic_vector(to_unsigned( 2840, 16)), --  2840 / 0x0b18
    5944 => std_logic_vector(to_unsigned( 4310, 16)), --  4310 / 0x10d6
    5945 => std_logic_vector(to_unsigned(  771, 16)), --   771 / 0x0303 -- last item of row
    5946 => std_logic_vector(to_unsigned( 4951, 16)), --  4951 / 0x1357
    5947 => std_logic_vector(to_unsigned(  211, 16)), --   211 / 0x00d3
    5948 => std_logic_vector(to_unsigned( 2208, 16)), --  2208 / 0x08a0
    5949 => std_logic_vector(to_unsigned(  723, 16)), --   723 / 0x02d3
    5950 => std_logic_vector(to_unsigned( 1246, 16)), --  1246 / 0x04de
    5951 => std_logic_vector(to_unsigned( 2928, 16)), --  2928 / 0x0b70
    5952 => std_logic_vector(to_unsigned(  398, 16)), --   398 / 0x018e
    5953 => std_logic_vector(to_unsigned( 5739, 16)), --  5739 / 0x166b
    5954 => std_logic_vector(to_unsigned(  265, 16)), --   265 / 0x0109
    5955 => std_logic_vector(to_unsigned( 5601, 16)), --  5601 / 0x15e1
    5956 => std_logic_vector(to_unsigned( 5993, 16)), --  5993 / 0x1769
    5957 => std_logic_vector(to_unsigned( 2615, 16)), --  2615 / 0x0a37 -- last item of row
    5958 => std_logic_vector(to_unsigned(  210, 16)), --   210 / 0x00d2
    5959 => std_logic_vector(to_unsigned( 4730, 16)), --  4730 / 0x127a
    5960 => std_logic_vector(to_unsigned( 5777, 16)), --  5777 / 0x1691
    5961 => std_logic_vector(to_unsigned( 3096, 16)), --  3096 / 0x0c18
    5962 => std_logic_vector(to_unsigned( 4282, 16)), --  4282 / 0x10ba
    5963 => std_logic_vector(to_unsigned( 6238, 16)), --  6238 / 0x185e
    5964 => std_logic_vector(to_unsigned( 4939, 16)), --  4939 / 0x134b
    5965 => std_logic_vector(to_unsigned( 1119, 16)), --  1119 / 0x045f
    5966 => std_logic_vector(to_unsigned( 6463, 16)), --  6463 / 0x193f
    5967 => std_logic_vector(to_unsigned( 5298, 16)), --  5298 / 0x14b2
    5968 => std_logic_vector(to_unsigned( 6320, 16)), --  6320 / 0x18b0
    5969 => std_logic_vector(to_unsigned( 4016, 16)), --  4016 / 0x0fb0 -- last item of row
    5970 => std_logic_vector(to_unsigned( 4167, 16)), --  4167 / 0x1047
    5971 => std_logic_vector(to_unsigned( 2063, 16)), --  2063 / 0x080f
    5972 => std_logic_vector(to_unsigned( 4757, 16)), --  4757 / 0x1295
    5973 => std_logic_vector(to_unsigned( 3157, 16)), --  3157 / 0x0c55
    5974 => std_logic_vector(to_unsigned( 5664, 16)), --  5664 / 0x1620
    5975 => std_logic_vector(to_unsigned( 3956, 16)), --  3956 / 0x0f74
    5976 => std_logic_vector(to_unsigned( 6045, 16)), --  6045 / 0x179d
    5977 => std_logic_vector(to_unsigned(  563, 16)), --   563 / 0x0233
    5978 => std_logic_vector(to_unsigned( 4284, 16)), --  4284 / 0x10bc
    5979 => std_logic_vector(to_unsigned( 2441, 16)), --  2441 / 0x0989
    5980 => std_logic_vector(to_unsigned( 3412, 16)), --  3412 / 0x0d54
    5981 => std_logic_vector(to_unsigned( 6334, 16)), --  6334 / 0x18be -- last item of row
    5982 => std_logic_vector(to_unsigned( 4201, 16)), --  4201 / 0x1069
    5983 => std_logic_vector(to_unsigned( 2428, 16)), --  2428 / 0x097c
    5984 => std_logic_vector(to_unsigned( 4474, 16)), --  4474 / 0x117a
    5985 => std_logic_vector(to_unsigned(   59, 16)), --    59 / 0x003b
    5986 => std_logic_vector(to_unsigned( 1721, 16)), --  1721 / 0x06b9
    5987 => std_logic_vector(to_unsigned(  736, 16)), --   736 / 0x02e0
    5988 => std_logic_vector(to_unsigned( 2997, 16)), --  2997 / 0x0bb5
    5989 => std_logic_vector(to_unsigned(  428, 16)), --   428 / 0x01ac
    5990 => std_logic_vector(to_unsigned( 3807, 16)), --  3807 / 0x0edf
    5991 => std_logic_vector(to_unsigned( 1513, 16)), --  1513 / 0x05e9
    5992 => std_logic_vector(to_unsigned( 4732, 16)), --  4732 / 0x127c
    5993 => std_logic_vector(to_unsigned( 6195, 16)), --  6195 / 0x1833 -- last item of row
    5994 => std_logic_vector(to_unsigned( 2670, 16)), --  2670 / 0x0a6e
    5995 => std_logic_vector(to_unsigned( 3081, 16)), --  3081 / 0x0c09
    5996 => std_logic_vector(to_unsigned( 5139, 16)), --  5139 / 0x1413
    5997 => std_logic_vector(to_unsigned( 3736, 16)), --  3736 / 0x0e98
    5998 => std_logic_vector(to_unsigned( 1999, 16)), --  1999 / 0x07cf
    5999 => std_logic_vector(to_unsigned( 5889, 16)), --  5889 / 0x1701
    6000 => std_logic_vector(to_unsigned( 4362, 16)), --  4362 / 0x110a
    6001 => std_logic_vector(to_unsigned( 3806, 16)), --  3806 / 0x0ede
    6002 => std_logic_vector(to_unsigned( 4534, 16)), --  4534 / 0x11b6
    6003 => std_logic_vector(to_unsigned( 5409, 16)), --  5409 / 0x1521
    6004 => std_logic_vector(to_unsigned( 6384, 16)), --  6384 / 0x18f0
    6005 => std_logic_vector(to_unsigned( 5809, 16)), --  5809 / 0x16b1 -- last item of row
    6006 => std_logic_vector(to_unsigned( 5516, 16)), --  5516 / 0x158c
    6007 => std_logic_vector(to_unsigned( 1622, 16)), --  1622 / 0x0656
    6008 => std_logic_vector(to_unsigned( 2906, 16)), --  2906 / 0x0b5a
    6009 => std_logic_vector(to_unsigned( 3285, 16)), --  3285 / 0x0cd5
    6010 => std_logic_vector(to_unsigned( 1257, 16)), --  1257 / 0x04e9
    6011 => std_logic_vector(to_unsigned( 5797, 16)), --  5797 / 0x16a5
    6012 => std_logic_vector(to_unsigned( 3816, 16)), --  3816 / 0x0ee8
    6013 => std_logic_vector(to_unsigned(  817, 16)), --   817 / 0x0331
    6014 => std_logic_vector(to_unsigned(  875, 16)), --   875 / 0x036b
    6015 => std_logic_vector(to_unsigned( 2311, 16)), --  2311 / 0x0907
    6016 => std_logic_vector(to_unsigned( 3543, 16)), --  3543 / 0x0dd7
    6017 => std_logic_vector(to_unsigned( 1205, 16)), --  1205 / 0x04b5 -- last item of row
    6018 => std_logic_vector(to_unsigned( 4244, 16)), --  4244 / 0x1094
    6019 => std_logic_vector(to_unsigned( 2184, 16)), --  2184 / 0x0888
    6020 => std_logic_vector(to_unsigned( 5415, 16)), --  5415 / 0x1527
    6021 => std_logic_vector(to_unsigned( 1705, 16)), --  1705 / 0x06a9
    6022 => std_logic_vector(to_unsigned( 5642, 16)), --  5642 / 0x160a
    6023 => std_logic_vector(to_unsigned( 4886, 16)), --  4886 / 0x1316
    6024 => std_logic_vector(to_unsigned( 2333, 16)), --  2333 / 0x091d
    6025 => std_logic_vector(to_unsigned(  287, 16)), --   287 / 0x011f
    6026 => std_logic_vector(to_unsigned( 1848, 16)), --  1848 / 0x0738
    6027 => std_logic_vector(to_unsigned( 1121, 16)), --  1121 / 0x0461
    6028 => std_logic_vector(to_unsigned( 3595, 16)), --  3595 / 0x0e0b
    6029 => std_logic_vector(to_unsigned( 6022, 16)), --  6022 / 0x1786 -- last item of row
    6030 => std_logic_vector(to_unsigned( 2142, 16)), --  2142 / 0x085e
    6031 => std_logic_vector(to_unsigned( 2830, 16)), --  2830 / 0x0b0e
    6032 => std_logic_vector(to_unsigned( 4069, 16)), --  4069 / 0x0fe5
    6033 => std_logic_vector(to_unsigned( 5654, 16)), --  5654 / 0x1616
    6034 => std_logic_vector(to_unsigned( 1295, 16)), --  1295 / 0x050f
    6035 => std_logic_vector(to_unsigned( 2951, 16)), --  2951 / 0x0b87
    6036 => std_logic_vector(to_unsigned( 3919, 16)), --  3919 / 0x0f4f
    6037 => std_logic_vector(to_unsigned( 1356, 16)), --  1356 / 0x054c
    6038 => std_logic_vector(to_unsigned(  884, 16)), --   884 / 0x0374
    6039 => std_logic_vector(to_unsigned( 1786, 16)), --  1786 / 0x06fa
    6040 => std_logic_vector(to_unsigned(  396, 16)), --   396 / 0x018c
    6041 => std_logic_vector(to_unsigned( 4738, 16)), --  4738 / 0x1282 -- last item of row
    6042 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6043 => std_logic_vector(to_unsigned( 2161, 16)), --  2161 / 0x0871
    6044 => std_logic_vector(to_unsigned( 2653, 16)), --  2653 / 0x0a5d -- last item of row
    6045 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6046 => std_logic_vector(to_unsigned( 1380, 16)), --  1380 / 0x0564
    6047 => std_logic_vector(to_unsigned( 1461, 16)), --  1461 / 0x05b5 -- last item of row
    6048 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6049 => std_logic_vector(to_unsigned( 2502, 16)), --  2502 / 0x09c6
    6050 => std_logic_vector(to_unsigned( 3707, 16)), --  3707 / 0x0e7b -- last item of row
    6051 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6052 => std_logic_vector(to_unsigned( 3971, 16)), --  3971 / 0x0f83
    6053 => std_logic_vector(to_unsigned( 1057, 16)), --  1057 / 0x0421 -- last item of row
    6054 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6055 => std_logic_vector(to_unsigned( 5985, 16)), --  5985 / 0x1761
    6056 => std_logic_vector(to_unsigned( 6062, 16)), --  6062 / 0x17ae -- last item of row
    6057 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6058 => std_logic_vector(to_unsigned( 1733, 16)), --  1733 / 0x06c5
    6059 => std_logic_vector(to_unsigned( 6028, 16)), --  6028 / 0x178c -- last item of row
    6060 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6061 => std_logic_vector(to_unsigned( 3786, 16)), --  3786 / 0x0eca
    6062 => std_logic_vector(to_unsigned( 1936, 16)), --  1936 / 0x0790 -- last item of row
    6063 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6064 => std_logic_vector(to_unsigned( 4292, 16)), --  4292 / 0x10c4
    6065 => std_logic_vector(to_unsigned(  956, 16)), --   956 / 0x03bc -- last item of row
    6066 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    6067 => std_logic_vector(to_unsigned( 5692, 16)), --  5692 / 0x163c
    6068 => std_logic_vector(to_unsigned( 3417, 16)), --  3417 / 0x0d59 -- last item of row
    6069 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    6070 => std_logic_vector(to_unsigned(  266, 16)), --   266 / 0x010a
    6071 => std_logic_vector(to_unsigned( 4878, 16)), --  4878 / 0x130e -- last item of row
    6072 => std_logic_vector(to_unsigned(   10, 16)), --    10 / 0x000a
    6073 => std_logic_vector(to_unsigned( 4913, 16)), --  4913 / 0x1331
    6074 => std_logic_vector(to_unsigned( 3247, 16)), --  3247 / 0x0caf -- last item of row
    6075 => std_logic_vector(to_unsigned(   11, 16)), --    11 / 0x000b
    6076 => std_logic_vector(to_unsigned( 4763, 16)), --  4763 / 0x129b
    6077 => std_logic_vector(to_unsigned( 3937, 16)), --  3937 / 0x0f61 -- last item of row
    6078 => std_logic_vector(to_unsigned(   12, 16)), --    12 / 0x000c
    6079 => std_logic_vector(to_unsigned( 3590, 16)), --  3590 / 0x0e06
    6080 => std_logic_vector(to_unsigned( 2903, 16)), --  2903 / 0x0b57 -- last item of row
    6081 => std_logic_vector(to_unsigned(   13, 16)), --    13 / 0x000d
    6082 => std_logic_vector(to_unsigned( 2566, 16)), --  2566 / 0x0a06
    6083 => std_logic_vector(to_unsigned( 4215, 16)), --  4215 / 0x1077 -- last item of row
    6084 => std_logic_vector(to_unsigned(   14, 16)), --    14 / 0x000e
    6085 => std_logic_vector(to_unsigned( 5208, 16)), --  5208 / 0x1458
    6086 => std_logic_vector(to_unsigned( 4707, 16)), --  4707 / 0x1263 -- last item of row
    6087 => std_logic_vector(to_unsigned(   15, 16)), --    15 / 0x000f
    6088 => std_logic_vector(to_unsigned( 3940, 16)), --  3940 / 0x0f64
    6089 => std_logic_vector(to_unsigned( 3388, 16)), --  3388 / 0x0d3c -- last item of row
    6090 => std_logic_vector(to_unsigned(   16, 16)), --    16 / 0x0010
    6091 => std_logic_vector(to_unsigned( 5109, 16)), --  5109 / 0x13f5
    6092 => std_logic_vector(to_unsigned( 4556, 16)), --  4556 / 0x11cc -- last item of row
    6093 => std_logic_vector(to_unsigned(   17, 16)), --    17 / 0x0011
    6094 => std_logic_vector(to_unsigned( 4908, 16)), --  4908 / 0x132c
    6095 => std_logic_vector(to_unsigned( 4177, 16)), --  4177 / 0x1051 -- last item of row
    -- Table for fecframe_short, C4_5
    6096 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6097 => std_logic_vector(to_unsigned(  896, 16)), --   896 / 0x0380
    6098 => std_logic_vector(to_unsigned( 1565, 16)), --  1565 / 0x061d -- last item of row
    6099 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6100 => std_logic_vector(to_unsigned( 2493, 16)), --  2493 / 0x09bd
    6101 => std_logic_vector(to_unsigned(  184, 16)), --   184 / 0x00b8 -- last item of row
    6102 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6103 => std_logic_vector(to_unsigned(  212, 16)), --   212 / 0x00d4
    6104 => std_logic_vector(to_unsigned( 3210, 16)), --  3210 / 0x0c8a -- last item of row
    6105 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    6106 => std_logic_vector(to_unsigned(  727, 16)), --   727 / 0x02d7
    6107 => std_logic_vector(to_unsigned( 1339, 16)), --  1339 / 0x053b -- last item of row
    6108 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    6109 => std_logic_vector(to_unsigned( 3428, 16)), --  3428 / 0x0d64
    6110 => std_logic_vector(to_unsigned(  612, 16)), --   612 / 0x0264 -- last item of row
    6111 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6112 => std_logic_vector(to_unsigned( 2663, 16)), --  2663 / 0x0a67
    6113 => std_logic_vector(to_unsigned( 1947, 16)), --  1947 / 0x079b -- last item of row
    6114 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6115 => std_logic_vector(to_unsigned(  230, 16)), --   230 / 0x00e6
    6116 => std_logic_vector(to_unsigned( 2695, 16)), --  2695 / 0x0a87 -- last item of row
    6117 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6118 => std_logic_vector(to_unsigned( 2025, 16)), --  2025 / 0x07e9
    6119 => std_logic_vector(to_unsigned( 2794, 16)), --  2794 / 0x0aea -- last item of row
    6120 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6121 => std_logic_vector(to_unsigned( 3039, 16)), --  3039 / 0x0bdf
    6122 => std_logic_vector(to_unsigned(  283, 16)), --   283 / 0x011b -- last item of row
    6123 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6124 => std_logic_vector(to_unsigned(  862, 16)), --   862 / 0x035e
    6125 => std_logic_vector(to_unsigned( 2889, 16)), --  2889 / 0x0b49 -- last item of row
    6126 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6127 => std_logic_vector(to_unsigned(  376, 16)), --   376 / 0x0178
    6128 => std_logic_vector(to_unsigned( 2110, 16)), --  2110 / 0x083e -- last item of row
    6129 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6130 => std_logic_vector(to_unsigned( 2034, 16)), --  2034 / 0x07f2
    6131 => std_logic_vector(to_unsigned( 2286, 16)), --  2286 / 0x08ee -- last item of row
    6132 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6133 => std_logic_vector(to_unsigned(  951, 16)), --   951 / 0x03b7
    6134 => std_logic_vector(to_unsigned( 2068, 16)), --  2068 / 0x0814 -- last item of row
    6135 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    6136 => std_logic_vector(to_unsigned( 3108, 16)), --  3108 / 0x0c24
    6137 => std_logic_vector(to_unsigned( 3542, 16)), --  3542 / 0x0dd6 -- last item of row
    6138 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    6139 => std_logic_vector(to_unsigned(  307, 16)), --   307 / 0x0133
    6140 => std_logic_vector(to_unsigned( 1421, 16)), --  1421 / 0x058d -- last item of row
    6141 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6142 => std_logic_vector(to_unsigned( 2272, 16)), --  2272 / 0x08e0
    6143 => std_logic_vector(to_unsigned( 1197, 16)), --  1197 / 0x04ad -- last item of row
    6144 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6145 => std_logic_vector(to_unsigned( 1800, 16)), --  1800 / 0x0708
    6146 => std_logic_vector(to_unsigned( 3280, 16)), --  3280 / 0x0cd0 -- last item of row
    6147 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6148 => std_logic_vector(to_unsigned(  331, 16)), --   331 / 0x014b
    6149 => std_logic_vector(to_unsigned( 2308, 16)), --  2308 / 0x0904 -- last item of row
    6150 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6151 => std_logic_vector(to_unsigned(  465, 16)), --   465 / 0x01d1
    6152 => std_logic_vector(to_unsigned( 2552, 16)), --  2552 / 0x09f8 -- last item of row
    6153 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6154 => std_logic_vector(to_unsigned( 1038, 16)), --  1038 / 0x040e
    6155 => std_logic_vector(to_unsigned( 2479, 16)), --  2479 / 0x09af -- last item of row
    6156 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6157 => std_logic_vector(to_unsigned( 1383, 16)), --  1383 / 0x0567
    6158 => std_logic_vector(to_unsigned(  343, 16)), --   343 / 0x0157 -- last item of row
    6159 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6160 => std_logic_vector(to_unsigned(   94, 16)), --    94 / 0x005e
    6161 => std_logic_vector(to_unsigned(  236, 16)), --   236 / 0x00ec -- last item of row
    6162 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6163 => std_logic_vector(to_unsigned( 2619, 16)), --  2619 / 0x0a3b
    6164 => std_logic_vector(to_unsigned(  121, 16)), --   121 / 0x0079 -- last item of row
    6165 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    6166 => std_logic_vector(to_unsigned( 1497, 16)), --  1497 / 0x05d9
    6167 => std_logic_vector(to_unsigned( 2774, 16)), --  2774 / 0x0ad6 -- last item of row
    6168 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    6169 => std_logic_vector(to_unsigned( 2116, 16)), --  2116 / 0x0844
    6170 => std_logic_vector(to_unsigned( 1855, 16)), --  1855 / 0x073f -- last item of row
    6171 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6172 => std_logic_vector(to_unsigned(  722, 16)), --   722 / 0x02d2
    6173 => std_logic_vector(to_unsigned( 1584, 16)), --  1584 / 0x0630 -- last item of row
    6174 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6175 => std_logic_vector(to_unsigned( 2767, 16)), --  2767 / 0x0acf
    6176 => std_logic_vector(to_unsigned( 1881, 16)), --  1881 / 0x0759 -- last item of row
    6177 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6178 => std_logic_vector(to_unsigned( 2701, 16)), --  2701 / 0x0a8d
    6179 => std_logic_vector(to_unsigned( 1610, 16)), --  1610 / 0x064a -- last item of row
    6180 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6181 => std_logic_vector(to_unsigned( 3283, 16)), --  3283 / 0x0cd3
    6182 => std_logic_vector(to_unsigned( 1732, 16)), --  1732 / 0x06c4 -- last item of row
    6183 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6184 => std_logic_vector(to_unsigned(  168, 16)), --   168 / 0x00a8
    6185 => std_logic_vector(to_unsigned( 1099, 16)), --  1099 / 0x044b -- last item of row
    6186 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6187 => std_logic_vector(to_unsigned( 3074, 16)), --  3074 / 0x0c02
    6188 => std_logic_vector(to_unsigned(  243, 16)), --   243 / 0x00f3 -- last item of row
    6189 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6190 => std_logic_vector(to_unsigned( 3460, 16)), --  3460 / 0x0d84
    6191 => std_logic_vector(to_unsigned(  945, 16)), --   945 / 0x03b1 -- last item of row
    6192 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6193 => std_logic_vector(to_unsigned( 2049, 16)), --  2049 / 0x0801
    6194 => std_logic_vector(to_unsigned( 1746, 16)), --  1746 / 0x06d2 -- last item of row
    6195 => std_logic_vector(to_unsigned(    8, 16)), --     8 / 0x0008
    6196 => std_logic_vector(to_unsigned(  566, 16)), --   566 / 0x0236
    6197 => std_logic_vector(to_unsigned( 1427, 16)), --  1427 / 0x0593 -- last item of row
    6198 => std_logic_vector(to_unsigned(    9, 16)), --     9 / 0x0009
    6199 => std_logic_vector(to_unsigned( 3545, 16)), --  3545 / 0x0dd9
    6200 => std_logic_vector(to_unsigned( 1168, 16)), --  1168 / 0x0490 -- last item of row
    -- Table for fecframe_short, C5_6
    6201 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6202 => std_logic_vector(to_unsigned( 2409, 16)), --  2409 / 0x0969
    6203 => std_logic_vector(to_unsigned(  499, 16)), --   499 / 0x01f3
    6204 => std_logic_vector(to_unsigned( 1481, 16)), --  1481 / 0x05c9
    6205 => std_logic_vector(to_unsigned(  908, 16)), --   908 / 0x038c
    6206 => std_logic_vector(to_unsigned(  559, 16)), --   559 / 0x022f
    6207 => std_logic_vector(to_unsigned(  716, 16)), --   716 / 0x02cc
    6208 => std_logic_vector(to_unsigned( 1270, 16)), --  1270 / 0x04f6
    6209 => std_logic_vector(to_unsigned(  333, 16)), --   333 / 0x014d
    6210 => std_logic_vector(to_unsigned( 2508, 16)), --  2508 / 0x09cc
    6211 => std_logic_vector(to_unsigned( 2264, 16)), --  2264 / 0x08d8
    6212 => std_logic_vector(to_unsigned( 1702, 16)), --  1702 / 0x06a6
    6213 => std_logic_vector(to_unsigned( 2805, 16)), --  2805 / 0x0af5 -- last item of row
    6214 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6215 => std_logic_vector(to_unsigned( 2447, 16)), --  2447 / 0x098f
    6216 => std_logic_vector(to_unsigned( 1926, 16)), --  1926 / 0x0786 -- last item of row
    6217 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6218 => std_logic_vector(to_unsigned(  414, 16)), --   414 / 0x019e
    6219 => std_logic_vector(to_unsigned( 1224, 16)), --  1224 / 0x04c8 -- last item of row
    6220 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6221 => std_logic_vector(to_unsigned( 2114, 16)), --  2114 / 0x0842
    6222 => std_logic_vector(to_unsigned(  842, 16)), --   842 / 0x034a -- last item of row
    6223 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6224 => std_logic_vector(to_unsigned(  212, 16)), --   212 / 0x00d4
    6225 => std_logic_vector(to_unsigned(  573, 16)), --   573 / 0x023d -- last item of row
    6226 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6227 => std_logic_vector(to_unsigned( 2383, 16)), --  2383 / 0x094f
    6228 => std_logic_vector(to_unsigned( 2112, 16)), --  2112 / 0x0840 -- last item of row
    6229 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6230 => std_logic_vector(to_unsigned( 2286, 16)), --  2286 / 0x08ee
    6231 => std_logic_vector(to_unsigned( 2348, 16)), --  2348 / 0x092c -- last item of row
    6232 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6233 => std_logic_vector(to_unsigned(  545, 16)), --   545 / 0x0221
    6234 => std_logic_vector(to_unsigned(  819, 16)), --   819 / 0x0333 -- last item of row
    6235 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6236 => std_logic_vector(to_unsigned( 1264, 16)), --  1264 / 0x04f0
    6237 => std_logic_vector(to_unsigned(  143, 16)), --   143 / 0x008f -- last item of row
    6238 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6239 => std_logic_vector(to_unsigned( 1701, 16)), --  1701 / 0x06a5
    6240 => std_logic_vector(to_unsigned( 2258, 16)), --  2258 / 0x08d2 -- last item of row
    6241 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6242 => std_logic_vector(to_unsigned(  964, 16)), --   964 / 0x03c4
    6243 => std_logic_vector(to_unsigned(  166, 16)), --   166 / 0x00a6 -- last item of row
    6244 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6245 => std_logic_vector(to_unsigned(  114, 16)), --   114 / 0x0072
    6246 => std_logic_vector(to_unsigned( 2413, 16)), --  2413 / 0x096d -- last item of row
    6247 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6248 => std_logic_vector(to_unsigned( 2243, 16)), --  2243 / 0x08c3
    6249 => std_logic_vector(to_unsigned(   81, 16)), --    81 / 0x0051 -- last item of row
    6250 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6251 => std_logic_vector(to_unsigned( 1245, 16)), --  1245 / 0x04dd
    6252 => std_logic_vector(to_unsigned( 1581, 16)), --  1581 / 0x062d -- last item of row
    6253 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6254 => std_logic_vector(to_unsigned(  775, 16)), --   775 / 0x0307
    6255 => std_logic_vector(to_unsigned(  169, 16)), --   169 / 0x00a9 -- last item of row
    6256 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6257 => std_logic_vector(to_unsigned( 1696, 16)), --  1696 / 0x06a0
    6258 => std_logic_vector(to_unsigned( 1104, 16)), --  1104 / 0x0450 -- last item of row
    6259 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6260 => std_logic_vector(to_unsigned( 1914, 16)), --  1914 / 0x077a
    6261 => std_logic_vector(to_unsigned( 2831, 16)), --  2831 / 0x0b0f -- last item of row
    6262 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6263 => std_logic_vector(to_unsigned(  532, 16)), --   532 / 0x0214
    6264 => std_logic_vector(to_unsigned( 1450, 16)), --  1450 / 0x05aa -- last item of row
    6265 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6266 => std_logic_vector(to_unsigned(   91, 16)), --    91 / 0x005b
    6267 => std_logic_vector(to_unsigned(  974, 16)), --   974 / 0x03ce -- last item of row
    6268 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6269 => std_logic_vector(to_unsigned(  497, 16)), --   497 / 0x01f1
    6270 => std_logic_vector(to_unsigned( 2228, 16)), --  2228 / 0x08b4 -- last item of row
    6271 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6272 => std_logic_vector(to_unsigned( 2326, 16)), --  2326 / 0x0916
    6273 => std_logic_vector(to_unsigned( 1579, 16)), --  1579 / 0x062b -- last item of row
    6274 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6275 => std_logic_vector(to_unsigned( 2482, 16)), --  2482 / 0x09b2
    6276 => std_logic_vector(to_unsigned(  256, 16)), --   256 / 0x0100 -- last item of row
    6277 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6278 => std_logic_vector(to_unsigned( 1117, 16)), --  1117 / 0x045d
    6279 => std_logic_vector(to_unsigned( 1261, 16)), --  1261 / 0x04ed -- last item of row
    6280 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6281 => std_logic_vector(to_unsigned( 1257, 16)), --  1257 / 0x04e9
    6282 => std_logic_vector(to_unsigned( 1658, 16)), --  1658 / 0x067a -- last item of row
    6283 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6284 => std_logic_vector(to_unsigned( 1478, 16)), --  1478 / 0x05c6
    6285 => std_logic_vector(to_unsigned( 1225, 16)), --  1225 / 0x04c9 -- last item of row
    6286 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6287 => std_logic_vector(to_unsigned( 2511, 16)), --  2511 / 0x09cf
    6288 => std_logic_vector(to_unsigned(  980, 16)), --   980 / 0x03d4 -- last item of row
    6289 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6290 => std_logic_vector(to_unsigned( 2320, 16)), --  2320 / 0x0910
    6291 => std_logic_vector(to_unsigned( 2675, 16)), --  2675 / 0x0a73 -- last item of row
    6292 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6293 => std_logic_vector(to_unsigned(  435, 16)), --   435 / 0x01b3
    6294 => std_logic_vector(to_unsigned( 1278, 16)), --  1278 / 0x04fe -- last item of row
    6295 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6296 => std_logic_vector(to_unsigned(  228, 16)), --   228 / 0x00e4
    6297 => std_logic_vector(to_unsigned(  503, 16)), --   503 / 0x01f7 -- last item of row
    6298 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6299 => std_logic_vector(to_unsigned( 1885, 16)), --  1885 / 0x075d
    6300 => std_logic_vector(to_unsigned( 2369, 16)), --  2369 / 0x0941 -- last item of row
    6301 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6302 => std_logic_vector(to_unsigned(   57, 16)), --    57 / 0x0039
    6303 => std_logic_vector(to_unsigned(  483, 16)), --   483 / 0x01e3 -- last item of row
    6304 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6305 => std_logic_vector(to_unsigned(  838, 16)), --   838 / 0x0346
    6306 => std_logic_vector(to_unsigned( 1050, 16)), --  1050 / 0x041a -- last item of row
    6307 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6308 => std_logic_vector(to_unsigned( 1231, 16)), --  1231 / 0x04cf
    6309 => std_logic_vector(to_unsigned( 1990, 16)), --  1990 / 0x07c6 -- last item of row
    6310 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6311 => std_logic_vector(to_unsigned( 1738, 16)), --  1738 / 0x06ca
    6312 => std_logic_vector(to_unsigned(   68, 16)), --    68 / 0x0044 -- last item of row
    6313 => std_logic_vector(to_unsigned(    5, 16)), --     5 / 0x0005
    6314 => std_logic_vector(to_unsigned( 2392, 16)), --  2392 / 0x0958
    6315 => std_logic_vector(to_unsigned(  951, 16)), --   951 / 0x03b7 -- last item of row
    6316 => std_logic_vector(to_unsigned(    6, 16)), --     6 / 0x0006
    6317 => std_logic_vector(to_unsigned(  163, 16)), --   163 / 0x00a3
    6318 => std_logic_vector(to_unsigned(  645, 16)), --   645 / 0x0285 -- last item of row
    6319 => std_logic_vector(to_unsigned(    7, 16)), --     7 / 0x0007
    6320 => std_logic_vector(to_unsigned( 2644, 16)), --  2644 / 0x0a54
    6321 => std_logic_vector(to_unsigned( 1704, 16)), --  1704 / 0x06a8 -- last item of row
    -- Table for fecframe_short, C8_9
    6322 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6323 => std_logic_vector(to_unsigned( 1558, 16)), --  1558 / 0x0616
    6324 => std_logic_vector(to_unsigned(  712, 16)), --   712 / 0x02c8
    6325 => std_logic_vector(to_unsigned(  805, 16)), --   805 / 0x0325 -- last item of row
    6326 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6327 => std_logic_vector(to_unsigned( 1450, 16)), --  1450 / 0x05aa
    6328 => std_logic_vector(to_unsigned(  873, 16)), --   873 / 0x0369
    6329 => std_logic_vector(to_unsigned( 1337, 16)), --  1337 / 0x0539 -- last item of row
    6330 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6331 => std_logic_vector(to_unsigned( 1741, 16)), --  1741 / 0x06cd
    6332 => std_logic_vector(to_unsigned( 1129, 16)), --  1129 / 0x0469
    6333 => std_logic_vector(to_unsigned( 1184, 16)), --  1184 / 0x04a0 -- last item of row
    6334 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6335 => std_logic_vector(to_unsigned(  294, 16)), --   294 / 0x0126
    6336 => std_logic_vector(to_unsigned(  806, 16)), --   806 / 0x0326
    6337 => std_logic_vector(to_unsigned( 1566, 16)), --  1566 / 0x061e -- last item of row
    6338 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6339 => std_logic_vector(to_unsigned(  482, 16)), --   482 / 0x01e2
    6340 => std_logic_vector(to_unsigned(  605, 16)), --   605 / 0x025d
    6341 => std_logic_vector(to_unsigned(  923, 16)), --   923 / 0x039b -- last item of row
    6342 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6343 => std_logic_vector(to_unsigned(  926, 16)), --   926 / 0x039e
    6344 => std_logic_vector(to_unsigned( 1578, 16)), --  1578 / 0x062a -- last item of row
    6345 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6346 => std_logic_vector(to_unsigned(  777, 16)), --   777 / 0x0309
    6347 => std_logic_vector(to_unsigned( 1374, 16)), --  1374 / 0x055e -- last item of row
    6348 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6349 => std_logic_vector(to_unsigned(  608, 16)), --   608 / 0x0260
    6350 => std_logic_vector(to_unsigned(  151, 16)), --   151 / 0x0097 -- last item of row
    6351 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6352 => std_logic_vector(to_unsigned( 1195, 16)), --  1195 / 0x04ab
    6353 => std_logic_vector(to_unsigned(  210, 16)), --   210 / 0x00d2 -- last item of row
    6354 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6355 => std_logic_vector(to_unsigned( 1484, 16)), --  1484 / 0x05cc
    6356 => std_logic_vector(to_unsigned(  692, 16)), --   692 / 0x02b4 -- last item of row
    6357 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6358 => std_logic_vector(to_unsigned(  427, 16)), --   427 / 0x01ab
    6359 => std_logic_vector(to_unsigned(  488, 16)), --   488 / 0x01e8 -- last item of row
    6360 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6361 => std_logic_vector(to_unsigned(  828, 16)), --   828 / 0x033c
    6362 => std_logic_vector(to_unsigned( 1124, 16)), --  1124 / 0x0464 -- last item of row
    6363 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6364 => std_logic_vector(to_unsigned(  874, 16)), --   874 / 0x036a
    6365 => std_logic_vector(to_unsigned( 1366, 16)), --  1366 / 0x0556 -- last item of row
    6366 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6367 => std_logic_vector(to_unsigned( 1500, 16)), --  1500 / 0x05dc
    6368 => std_logic_vector(to_unsigned(  835, 16)), --   835 / 0x0343 -- last item of row
    6369 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6370 => std_logic_vector(to_unsigned( 1496, 16)), --  1496 / 0x05d8
    6371 => std_logic_vector(to_unsigned(  502, 16)), --   502 / 0x01f6 -- last item of row
    6372 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6373 => std_logic_vector(to_unsigned( 1006, 16)), --  1006 / 0x03ee
    6374 => std_logic_vector(to_unsigned( 1701, 16)), --  1701 / 0x06a5 -- last item of row
    6375 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6376 => std_logic_vector(to_unsigned( 1155, 16)), --  1155 / 0x0483
    6377 => std_logic_vector(to_unsigned(   97, 16)), --    97 / 0x0061 -- last item of row
    6378 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6379 => std_logic_vector(to_unsigned(  657, 16)), --   657 / 0x0291
    6380 => std_logic_vector(to_unsigned( 1403, 16)), --  1403 / 0x057b -- last item of row
    6381 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6382 => std_logic_vector(to_unsigned( 1453, 16)), --  1453 / 0x05ad
    6383 => std_logic_vector(to_unsigned(  624, 16)), --   624 / 0x0270 -- last item of row
    6384 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6385 => std_logic_vector(to_unsigned(  429, 16)), --   429 / 0x01ad
    6386 => std_logic_vector(to_unsigned( 1495, 16)), --  1495 / 0x05d7 -- last item of row
    6387 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6388 => std_logic_vector(to_unsigned(  809, 16)), --   809 / 0x0329
    6389 => std_logic_vector(to_unsigned(  385, 16)), --   385 / 0x0181 -- last item of row
    6390 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6391 => std_logic_vector(to_unsigned(  367, 16)), --   367 / 0x016f
    6392 => std_logic_vector(to_unsigned(  151, 16)), --   151 / 0x0097 -- last item of row
    6393 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6394 => std_logic_vector(to_unsigned( 1323, 16)), --  1323 / 0x052b
    6395 => std_logic_vector(to_unsigned(  202, 16)), --   202 / 0x00ca -- last item of row
    6396 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6397 => std_logic_vector(to_unsigned(  960, 16)), --   960 / 0x03c0
    6398 => std_logic_vector(to_unsigned(  318, 16)), --   318 / 0x013e -- last item of row
    6399 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6400 => std_logic_vector(to_unsigned( 1451, 16)), --  1451 / 0x05ab
    6401 => std_logic_vector(to_unsigned( 1039, 16)), --  1039 / 0x040f -- last item of row
    6402 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6403 => std_logic_vector(to_unsigned( 1098, 16)), --  1098 / 0x044a
    6404 => std_logic_vector(to_unsigned( 1722, 16)), --  1722 / 0x06ba -- last item of row
    6405 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6406 => std_logic_vector(to_unsigned( 1015, 16)), --  1015 / 0x03f7
    6407 => std_logic_vector(to_unsigned( 1428, 16)), --  1428 / 0x0594 -- last item of row
    6408 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6409 => std_logic_vector(to_unsigned( 1261, 16)), --  1261 / 0x04ed
    6410 => std_logic_vector(to_unsigned( 1564, 16)), --  1564 / 0x061c -- last item of row
    6411 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6412 => std_logic_vector(to_unsigned(  544, 16)), --   544 / 0x0220
    6413 => std_logic_vector(to_unsigned( 1190, 16)), --  1190 / 0x04a6 -- last item of row
    6414 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6415 => std_logic_vector(to_unsigned( 1472, 16)), --  1472 / 0x05c0
    6416 => std_logic_vector(to_unsigned( 1246, 16)), --  1246 / 0x04de -- last item of row
    6417 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6418 => std_logic_vector(to_unsigned(  508, 16)), --   508 / 0x01fc
    6419 => std_logic_vector(to_unsigned(  630, 16)), --   630 / 0x0276 -- last item of row
    6420 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6421 => std_logic_vector(to_unsigned(  421, 16)), --   421 / 0x01a5
    6422 => std_logic_vector(to_unsigned( 1704, 16)), --  1704 / 0x06a8 -- last item of row
    6423 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6424 => std_logic_vector(to_unsigned(  284, 16)), --   284 / 0x011c
    6425 => std_logic_vector(to_unsigned(  898, 16)), --   898 / 0x0382 -- last item of row
    6426 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6427 => std_logic_vector(to_unsigned(  392, 16)), --   392 / 0x0188
    6428 => std_logic_vector(to_unsigned(  577, 16)), --   577 / 0x0241 -- last item of row
    6429 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6430 => std_logic_vector(to_unsigned( 1155, 16)), --  1155 / 0x0483
    6431 => std_logic_vector(to_unsigned(  556, 16)), --   556 / 0x022c -- last item of row
    6432 => std_logic_vector(to_unsigned(    0, 16)), --     0 / 0x0000
    6433 => std_logic_vector(to_unsigned(  631, 16)), --   631 / 0x0277
    6434 => std_logic_vector(to_unsigned( 1000, 16)), --  1000 / 0x03e8 -- last item of row
    6435 => std_logic_vector(to_unsigned(    1, 16)), --     1 / 0x0001
    6436 => std_logic_vector(to_unsigned(  732, 16)), --   732 / 0x02dc
    6437 => std_logic_vector(to_unsigned( 1368, 16)), --  1368 / 0x0558 -- last item of row
    6438 => std_logic_vector(to_unsigned(    2, 16)), --     2 / 0x0002
    6439 => std_logic_vector(to_unsigned( 1328, 16)), --  1328 / 0x0530
    6440 => std_logic_vector(to_unsigned(  329, 16)), --   329 / 0x0149 -- last item of row
    6441 => std_logic_vector(to_unsigned(    3, 16)), --     3 / 0x0003
    6442 => std_logic_vector(to_unsigned( 1515, 16)), --  1515 / 0x05eb
    6443 => std_logic_vector(to_unsigned(  506, 16)), --   506 / 0x01fa -- last item of row
    6444 => std_logic_vector(to_unsigned(    4, 16)), --     4 / 0x0004
    6445 => std_logic_vector(to_unsigned( 1104, 16)), --  1104 / 0x0450
    6446 => std_logic_vector(to_unsigned( 1172, 16)));

end package ldpc_tables_pkg;

package body ldpc_tables_pkg is
  -- Use this function to get the starting address of a given config within the LDPC_DATA_TABLE
  function get_ldpc_metadata (
    constant frame_length : frame_type_t;
    constant code_rate : code_rate_t) return ldpc_metadata_t is
  begin
    if frame_length = fecframe_normal and code_rate = C1_2 then
      return (
        addr => 0,
        q => 90,
        stage_0_loops => 36,
        stage_0_rows => 8,
        stage_1_loops => 54,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C1_3 then
      return (
        addr => 450,
        q => 120,
        stage_0_loops => 20,
        stage_0_rows => 12,
        stage_1_loops => 40,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C1_4 then
      return (
        addr => 810,
        q => 135,
        stage_0_loops => 15,
        stage_0_rows => 12,
        stage_1_loops => 30,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C2_3 then
      return (
        addr => 1080,
        q => 60,
        stage_0_loops => 12,
        stage_0_rows => 13,
        stage_1_loops => 108,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C2_5 then
      return (
        addr => 1560,
        q => 108,
        stage_0_loops => 24,
        stage_0_rows => 12,
        stage_1_loops => 48,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C3_4 then
      return (
        addr => 1992,
        q => 45,
        stage_0_loops => 15,
        stage_0_rows => 12,
        stage_1_loops => 120,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C3_5 then
      return (
        addr => 2532,
        q => 72,
        stage_0_loops => 36,
        stage_0_rows => 12,
        stage_1_loops => 72,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C4_5 then
      return (
        addr => 3180,
        q => 36,
        stage_0_loops => 18,
        stage_0_rows => 11,
        stage_1_loops => 126,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C5_6 then
      return (
        addr => 3756,
        q => 30,
        stage_0_loops => 15,
        stage_0_rows => 13,
        stage_1_loops => 135,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C8_9 then
      return (
        addr => 4356,
        q => 20,
        stage_0_loops => 20,
        stage_0_rows => 4,
        stage_1_loops => 140,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C9_10 then
      return (
        addr => 4856,
        q => 18,
        stage_0_loops => 18,
        stage_0_rows => 4,
        stage_1_loops => 144,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_2 then
      return (
        addr => 5360,
        q => 25,
        stage_0_loops => 5,
        stage_0_rows => 8,
        stage_1_loops => 15,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_3 then
      return (
        addr => 5445,
        q => 30,
        stage_0_loops => 5,
        stage_0_rows => 12,
        stage_1_loops => 10,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_4 then
      return (
        addr => 5535,
        q => 36,
        stage_0_loops => 4,
        stage_0_rows => 12,
        stage_1_loops => 5,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C2_3 then
      return (
        addr => 5598,
        q => 15,
        stage_0_loops => 3,
        stage_0_rows => 13,
        stage_1_loops => 27,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C2_5 then
      return (
        addr => 5718,
        q => 27,
        stage_0_loops => 6,
        stage_0_rows => 12,
        stage_1_loops => 12,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C3_4 then
      return (
        addr => 5826,
        q => 12,
        stage_0_loops => 1,
        stage_0_rows => 12,
        stage_1_loops => 32,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C3_5 then
      return (
        addr => 5934,
        q => 18,
        stage_0_loops => 9,
        stage_0_rows => 12,
        stage_1_loops => 18,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C4_5 then
      return (
        addr => 6096,
        q => 10,
        stage_0_loops => 17,
        stage_0_rows => 3,
        stage_1_loops => 18,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C5_6 then
      return (
        addr => 6201,
        q => 8,
        stage_0_loops => 1,
        stage_0_rows => 13,
        stage_1_loops => 36,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C8_9 then
      return (
        addr => 6322,
        q => 5,
        stage_0_loops => 5,
        stage_0_rows => 4,
        stage_1_loops => 35,
        stage_1_rows => 3);
     end if;

    -- Return a non existing index for any config not listed above
    return (addr => -1, q => -1, stage_0_loops => -1, stage_0_rows => -1, stage_1_loops => -1, stage_1_rows => -1);
  end function get_ldpc_metadata;

end package body ldpc_tables_pkg;