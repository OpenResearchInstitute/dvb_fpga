--    /*  -------------------------------------------------------------------------
--    This program is free software: you can redistribute it and/or modify
--    it under the terms of the GNU General Public License as published by
--    the Free Software Foundation, either version 3 of the License, or
--    any later version.
--
--    This program is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--    
--    You should have received a copy of the GNU General Public License
--    along with this program.  If not, see <http://www.gnu.org/licenses/>.
--    
--    Copyright: Levent Ozturk crc@leventozturk.com
--    https://leventozturk.com/engineering/crc/
--    Polynomial: x192+x190+x187+x186+x185+x181+x178+x177+x171+x170+x169+x167+x161+x160+x159+x154+x150+x148+x147+x146+x142+x140+x136+x132+x131+x130+x126+x124+x119+x118+x115+x114+x113+x112+x109+x107+x106+x103+x102+x100+x99+x95+x94+x92+x91+x90+x85+x84+x82+x80+x75+x71+x67+x64+x57+x56+x54+x50+x49+x48+x47+x42+x40+x39+x38+x37+x36+x34+x33+x32+x30+x29+x26+x25+x17+x14+x12+x10+x8+x7+x6+x5+x2+x1+1
--    d7 is the first data processed

--    c is internal LFSR state and the CRC output. Not needed for other modules than CRC.
--    c width is always same as polynomial width.
--    o is the output of all modules except CRC. Not needed for CRC.
--    o width is always same as data width width
-------------------------------------------------------------------------*/

-- Based on https://leventozturk.com/engineering/crc/

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bch_192x8 is generic (
	SEED : in std_ulogic_vector(191 downto 0) := (others => '0')
); port (
	clk   :  in std_ulogic;
	reset :  in std_ulogic;
	fd    :  in std_ulogic; -- First data. 1: SEED is used (initialise and calculate), 0: Previous CRC is used (continue and calculate)
	nd    :  in std_ulogic; -- New Data. d input has a valid data. Calculate new CRC
	rdy   : out std_ulogic;
	d    :  in std_ulogic_vector(  7 downto 0);  -- Data in
	c    : out std_ulogic_vector(191 downto 0);
 -- CRC output
    o    : out std_ulogic_vector(  7 downto 0) -- Data output
); end bch_192x8;

architecture a1 of bch_192x8 is
	signal                       nd_q : std_ulogic;
	signal                       fd_q : std_ulogic;
	signal                       dq : std_ulogic_vector (191 downto 0);
	signal                       ca : std_ulogic_vector(191 downto 0);
	signal                       oa : std_ulogic_vector(  7 downto 0);
begin
	process (clk)
	begin
		if (rising_edge(clk)) then
			nd_q <= nd;
			fd_q <= fd;
			dq(  0) <= d(  7) xor d(  5) xor d(  4) xor d(  2) xor d(  0);
			dq(  1) <= d(  7) xor d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(  2) <= d(  3) xor d(  1) xor d(  0);
			dq(  3) <= d(  4) xor d(  2) xor d(  1);
			dq(  4) <= d(  5) xor d(  3) xor d(  2);
			dq(  5) <= d(  7) xor d(  6) xor d(  5) xor d(  3) xor d(  2) xor d(  0);
			dq(  6) <= d(  6) xor d(  5) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(  7) <= d(  6) xor d(  5) xor d(  3) xor d(  1) xor d(  0);
			dq(  8) <= d(  6) xor d(  5) xor d(  1) xor d(  0);
			dq(  9) <= d(  7) xor d(  6) xor d(  2) xor d(  1);
			dq( 10) <= d(  5) xor d(  4) xor d(  3) xor d(  0);
			dq( 11) <= d(  6) xor d(  5) xor d(  4) xor d(  1);
			dq( 12) <= d(  6) xor d(  4) xor d(  0);
			dq( 13) <= d(  7) xor d(  5) xor d(  1);
			dq( 14) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  0);
			dq( 15) <= d(  7) xor d(  6) xor d(  5) xor d(  1);
			dq( 16) <= d(  7) xor d(  6) xor d(  2);
			dq( 17) <= d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  0);
			dq( 18) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  1);
			dq( 19) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  2);
			dq( 20) <= d(  7) xor d(  6) xor d(  5) xor d(  3);
			dq( 21) <= d(  7) xor d(  6) xor d(  4);
			dq( 22) <= d(  7) xor d(  5);
			dq( 23) <= d(  6);
			dq( 24) <= d(  7);
			dq( 25) <= d(  7) xor d(  5) xor d(  4) xor d(  2) xor d(  0);
			dq( 26) <= d(  7) xor d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq( 27) <= d(  7) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq( 28) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2);
			dq( 29) <= d(  6) xor d(  3) xor d(  2) xor d(  0);
			dq( 30) <= d(  5) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq( 31) <= d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq( 32) <= d(  3) xor d(  0);
			dq( 33) <= d(  7) xor d(  5) xor d(  2) xor d(  1) xor d(  0);
			dq( 34) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  1) xor d(  0);
			dq( 35) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  2) xor d(  1);
			dq( 36) <= d(  6) xor d(  4) xor d(  3) xor d(  0);
			dq( 37) <= d(  2) xor d(  1) xor d(  0);
			dq( 38) <= d(  7) xor d(  5) xor d(  4) xor d(  3) xor d(  1) xor d(  0);
			dq( 39) <= d(  7) xor d(  6) xor d(  1) xor d(  0);
			dq( 40) <= d(  5) xor d(  4) xor d(  1) xor d(  0);
			dq( 41) <= d(  6) xor d(  5) xor d(  2) xor d(  1);
			dq( 42) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  0);
			dq( 43) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  1);
			dq( 44) <= d(  7) xor d(  6) xor d(  5) xor d(  2);
			dq( 45) <= d(  7) xor d(  6) xor d(  3);
			dq( 46) <= d(  7) xor d(  4);
			dq( 47) <= d(  7) xor d(  4) xor d(  2) xor d(  0);
			dq( 48) <= d(  7) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq( 49) <= d(  7) xor d(  3) xor d(  1) xor d(  0);
			dq( 50) <= d(  7) xor d(  5) xor d(  1) xor d(  0);
			dq( 51) <= d(  6) xor d(  2) xor d(  1);
			dq( 52) <= d(  7) xor d(  3) xor d(  2);
			dq( 53) <= d(  4) xor d(  3);
			dq( 54) <= d(  7) xor d(  2) xor d(  0);
			dq( 55) <= d(  3) xor d(  1);
			dq( 56) <= d(  7) xor d(  5) xor d(  0);
			dq( 57) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  2) xor d(  1) xor d(  0);
			dq( 58) <= d(  7) xor d(  6) xor d(  5) xor d(  3) xor d(  2) xor d(  1);
			dq( 59) <= d(  7) xor d(  6) xor d(  4) xor d(  3) xor d(  2);
			dq( 60) <= d(  7) xor d(  5) xor d(  4) xor d(  3);
			dq( 61) <= d(  6) xor d(  5) xor d(  4);
			dq( 62) <= d(  7) xor d(  6) xor d(  5);
			dq( 63) <= d(  7) xor d(  6);
			dq( 64) <= d(  5) xor d(  4) xor d(  2) xor d(  0);
			dq( 65) <= d(  6) xor d(  5) xor d(  3) xor d(  1);
			dq( 66) <= d(  7) xor d(  6) xor d(  4) xor d(  2);
			dq( 67) <= d(  4) xor d(  3) xor d(  2) xor d(  0);
			dq( 68) <= d(  5) xor d(  4) xor d(  3) xor d(  1);
			dq( 69) <= d(  6) xor d(  5) xor d(  4) xor d(  2);
			dq( 70) <= d(  7) xor d(  6) xor d(  5) xor d(  3);
			dq( 71) <= d(  6) xor d(  5) xor d(  2) xor d(  0);
			dq( 72) <= d(  7) xor d(  6) xor d(  3) xor d(  1);
			dq( 73) <= d(  7) xor d(  4) xor d(  2);
			dq( 74) <= d(  5) xor d(  3);
			dq( 75) <= d(  7) xor d(  6) xor d(  5) xor d(  2) xor d(  0);
			dq( 76) <= d(  7) xor d(  6) xor d(  3) xor d(  1);
			dq( 77) <= d(  7) xor d(  4) xor d(  2);
			dq( 78) <= d(  5) xor d(  3);
			dq( 79) <= d(  6) xor d(  4);
			dq( 80) <= d(  4) xor d(  2) xor d(  0);
			dq( 81) <= d(  5) xor d(  3) xor d(  1);
			dq( 82) <= d(  7) xor d(  6) xor d(  5) xor d(  0);
			dq( 83) <= d(  7) xor d(  6) xor d(  1);
			dq( 84) <= d(  5) xor d(  4) xor d(  0);
			dq( 85) <= d(  7) xor d(  6) xor d(  4) xor d(  2) xor d(  1) xor d(  0);
			dq( 86) <= d(  7) xor d(  5) xor d(  3) xor d(  2) xor d(  1);
			dq( 87) <= d(  6) xor d(  4) xor d(  3) xor d(  2);
			dq( 88) <= d(  7) xor d(  5) xor d(  4) xor d(  3);
			dq( 89) <= d(  6) xor d(  5) xor d(  4);
			dq( 90) <= d(  6) xor d(  4) xor d(  2) xor d(  0);
			dq( 91) <= d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq( 92) <= d(  7) xor d(  3) xor d(  1) xor d(  0);
			dq( 93) <= d(  4) xor d(  2) xor d(  1);
			dq( 94) <= d(  7) xor d(  4) xor d(  3) xor d(  0);
			dq( 95) <= d(  7) xor d(  2) xor d(  1) xor d(  0);
			dq( 96) <= d(  3) xor d(  2) xor d(  1);
			dq( 97) <= d(  4) xor d(  3) xor d(  2);
			dq( 98) <= d(  5) xor d(  4) xor d(  3);
			dq( 99) <= d(  7) xor d(  6) xor d(  2) xor d(  0);
			dq(100) <= d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(101) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq(102) <= d(  6) xor d(  3) xor d(  0);
			dq(103) <= d(  5) xor d(  2) xor d(  1) xor d(  0);
			dq(104) <= d(  6) xor d(  3) xor d(  2) xor d(  1);
			dq(105) <= d(  7) xor d(  4) xor d(  3) xor d(  2);
			dq(106) <= d(  7) xor d(  3) xor d(  2) xor d(  0);
			dq(107) <= d(  7) xor d(  5) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(108) <= d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq(109) <= d(  3) xor d(  0);
			dq(110) <= d(  4) xor d(  1);
			dq(111) <= d(  5) xor d(  2);
			dq(112) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  0);
			dq(113) <= d(  6) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(114) <= d(  5) xor d(  3) xor d(  1) xor d(  0);
			dq(115) <= d(  7) xor d(  6) xor d(  5) xor d(  1) xor d(  0);
			dq(116) <= d(  7) xor d(  6) xor d(  2) xor d(  1);
			dq(117) <= d(  7) xor d(  3) xor d(  2);
			dq(118) <= d(  7) xor d(  5) xor d(  3) xor d(  2) xor d(  0);
			dq(119) <= d(  7) xor d(  6) xor d(  5) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(120) <= d(  7) xor d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq(121) <= d(  7) xor d(  5) xor d(  4) xor d(  3) xor d(  2);
			dq(122) <= d(  6) xor d(  5) xor d(  4) xor d(  3);
			dq(123) <= d(  7) xor d(  6) xor d(  5) xor d(  4);
			dq(124) <= d(  6) xor d(  4) xor d(  2) xor d(  0);
			dq(125) <= d(  7) xor d(  5) xor d(  3) xor d(  1);
			dq(126) <= d(  7) xor d(  6) xor d(  5) xor d(  0);
			dq(127) <= d(  7) xor d(  6) xor d(  1);
			dq(128) <= d(  7) xor d(  2);
			dq(129) <= d(  3);
			dq(130) <= d(  7) xor d(  5) xor d(  2) xor d(  0);
			dq(131) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(132) <= d(  6) xor d(  3) xor d(  1) xor d(  0);
			dq(133) <= d(  7) xor d(  4) xor d(  2) xor d(  1);
			dq(134) <= d(  5) xor d(  3) xor d(  2);
			dq(135) <= d(  6) xor d(  4) xor d(  3);
			dq(136) <= d(  2) xor d(  0);
			dq(137) <= d(  3) xor d(  1);
			dq(138) <= d(  4) xor d(  2);
			dq(139) <= d(  5) xor d(  3);
			dq(140) <= d(  7) xor d(  6) xor d(  5) xor d(  2) xor d(  0);
			dq(141) <= d(  7) xor d(  6) xor d(  3) xor d(  1);
			dq(142) <= d(  5) xor d(  0);
			dq(143) <= d(  6) xor d(  1);
			dq(144) <= d(  7) xor d(  2);
			dq(145) <= d(  3);
			dq(146) <= d(  7) xor d(  5) xor d(  2) xor d(  0);
			dq(147) <= d(  7) xor d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(148) <= d(  6) xor d(  3) xor d(  1) xor d(  0);
			dq(149) <= d(  7) xor d(  4) xor d(  2) xor d(  1);
			dq(150) <= d(  7) xor d(  4) xor d(  3) xor d(  0);
			dq(151) <= d(  5) xor d(  4) xor d(  1);
			dq(152) <= d(  6) xor d(  5) xor d(  2);
			dq(153) <= d(  7) xor d(  6) xor d(  3);
			dq(154) <= d(  5) xor d(  2) xor d(  0);
			dq(155) <= d(  6) xor d(  3) xor d(  1);
			dq(156) <= d(  7) xor d(  4) xor d(  2);
			dq(157) <= d(  5) xor d(  3);
			dq(158) <= d(  6) xor d(  4);
			dq(159) <= d(  4) xor d(  2) xor d(  0);
			dq(160) <= d(  7) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(161) <= d(  7) xor d(  3) xor d(  1) xor d(  0);
			dq(162) <= d(  4) xor d(  2) xor d(  1);
			dq(163) <= d(  5) xor d(  3) xor d(  2);
			dq(164) <= d(  6) xor d(  4) xor d(  3);
			dq(165) <= d(  7) xor d(  5) xor d(  4);
			dq(166) <= d(  6) xor d(  5);
			dq(167) <= d(  6) xor d(  5) xor d(  4) xor d(  2) xor d(  0);
			dq(168) <= d(  7) xor d(  6) xor d(  5) xor d(  3) xor d(  1);
			dq(169) <= d(  6) xor d(  5) xor d(  0);
			dq(170) <= d(  6) xor d(  5) xor d(  4) xor d(  2) xor d(  1) xor d(  0);
			dq(171) <= d(  6) xor d(  4) xor d(  3) xor d(  1) xor d(  0);
			dq(172) <= d(  7) xor d(  5) xor d(  4) xor d(  2) xor d(  1);
			dq(173) <= d(  6) xor d(  5) xor d(  3) xor d(  2);
			dq(174) <= d(  7) xor d(  6) xor d(  4) xor d(  3);
			dq(175) <= d(  7) xor d(  5) xor d(  4);
			dq(176) <= d(  6) xor d(  5);
			dq(177) <= d(  6) xor d(  5) xor d(  4) xor d(  2) xor d(  0);
			dq(178) <= d(  6) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(179) <= d(  7) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1);
			dq(180) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2);
			dq(181) <= d(  6) xor d(  3) xor d(  2) xor d(  0);
			dq(182) <= d(  7) xor d(  4) xor d(  3) xor d(  1);
			dq(183) <= d(  5) xor d(  4) xor d(  2);
			dq(184) <= d(  6) xor d(  5) xor d(  3);
			dq(185) <= d(  6) xor d(  5) xor d(  2) xor d(  0);
			dq(186) <= d(  6) xor d(  5) xor d(  4) xor d(  3) xor d(  2) xor d(  1) xor d(  0);
			dq(187) <= d(  6) xor d(  3) xor d(  1) xor d(  0);
			dq(188) <= d(  7) xor d(  4) xor d(  2) xor d(  1);
			dq(189) <= d(  5) xor d(  3) xor d(  2);
			dq(190) <= d(  7) xor d(  6) xor d(  5) xor d(  3) xor d(  2) xor d(  0);
			dq(191) <= d(  7) xor d(  6) xor d(  4) xor d(  3) xor d(  1);

		end if;
	end process;

	process (clk, reset)
	begin
		if (reset= '1') then
			ca <= SEED;
			rdy <= '0';
		elsif (rising_edge(clk)) then
			rdy <= nd_q;
			if(nd_q= '1') then
				if (fd_q= '1') then
					ca(  0) <= SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(  0);
					ca(  1) <= SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq(  1);
					ca(  2) <= SEED(184) xor SEED(185) xor SEED(187) xor dq(  2);
					ca(  3) <= SEED(185) xor SEED(186) xor SEED(188) xor dq(  3);
					ca(  4) <= SEED(186) xor SEED(187) xor SEED(189) xor dq(  4);
					ca(  5) <= SEED(184) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(  5);
					ca(  6) <= SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor dq(  6);
					ca(  7) <= SEED(184) xor SEED(185) xor SEED(187) xor SEED(189) xor SEED(190) xor dq(  7);
					ca(  8) <= SEED(  0) xor SEED(184) xor SEED(185) xor SEED(189) xor SEED(190) xor dq(  8);
					ca(  9) <= SEED(  1) xor SEED(185) xor SEED(186) xor SEED(190) xor SEED(191) xor dq(  9);
					ca( 10) <= SEED(  2) xor SEED(184) xor SEED(187) xor SEED(188) xor SEED(189) xor dq( 10);
					ca( 11) <= SEED(  3) xor SEED(185) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 11);
					ca( 12) <= SEED(  4) xor SEED(184) xor SEED(188) xor SEED(190) xor dq( 12);
					ca( 13) <= SEED(  5) xor SEED(185) xor SEED(189) xor SEED(191) xor dq( 13);
					ca( 14) <= SEED(  6) xor SEED(184) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 14);
					ca( 15) <= SEED(  7) xor SEED(185) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 15);
					ca( 16) <= SEED(  8) xor SEED(186) xor SEED(190) xor SEED(191) xor dq( 16);
					ca( 17) <= SEED(  9) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor dq( 17);
					ca( 18) <= SEED( 10) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 18);
					ca( 19) <= SEED( 11) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 19);
					ca( 20) <= SEED( 12) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 20);
					ca( 21) <= SEED( 13) xor SEED(188) xor SEED(190) xor SEED(191) xor dq( 21);
					ca( 22) <= SEED( 14) xor SEED(189) xor SEED(191) xor dq( 22);
					ca( 23) <= SEED( 15) xor SEED(190) xor dq( 23);
					ca( 24) <= SEED( 16) xor SEED(191) xor dq( 24);
					ca( 25) <= SEED( 17) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(191) xor dq( 25);
					ca( 26) <= SEED( 18) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq( 26);
					ca( 27) <= SEED( 19) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq( 27);
					ca( 28) <= SEED( 20) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 28);
					ca( 29) <= SEED( 21) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(190) xor dq( 29);
					ca( 30) <= SEED( 22) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor dq( 30);
					ca( 31) <= SEED( 23) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor dq( 31);
					ca( 32) <= SEED( 24) xor SEED(184) xor SEED(187) xor dq( 32);
					ca( 33) <= SEED( 25) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(189) xor SEED(191) xor dq( 33);
					ca( 34) <= SEED( 26) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 34);
					ca( 35) <= SEED( 27) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 35);
					ca( 36) <= SEED( 28) xor SEED(184) xor SEED(187) xor SEED(188) xor SEED(190) xor dq( 36);
					ca( 37) <= SEED( 29) xor SEED(184) xor SEED(185) xor SEED(186) xor dq( 37);
					ca( 38) <= SEED( 30) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq( 38);
					ca( 39) <= SEED( 31) xor SEED(184) xor SEED(185) xor SEED(190) xor SEED(191) xor dq( 39);
					ca( 40) <= SEED( 32) xor SEED(184) xor SEED(185) xor SEED(188) xor SEED(189) xor dq( 40);
					ca( 41) <= SEED( 33) xor SEED(185) xor SEED(186) xor SEED(189) xor SEED(190) xor dq( 41);
					ca( 42) <= SEED( 34) xor SEED(184) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 42);
					ca( 43) <= SEED( 35) xor SEED(185) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 43);
					ca( 44) <= SEED( 36) xor SEED(186) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 44);
					ca( 45) <= SEED( 37) xor SEED(187) xor SEED(190) xor SEED(191) xor dq( 45);
					ca( 46) <= SEED( 38) xor SEED(188) xor SEED(191) xor dq( 46);
					ca( 47) <= SEED( 39) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(191) xor dq( 47);
					ca( 48) <= SEED( 40) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(191) xor dq( 48);
					ca( 49) <= SEED( 41) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(191) xor dq( 49);
					ca( 50) <= SEED( 42) xor SEED(184) xor SEED(185) xor SEED(189) xor SEED(191) xor dq( 50);
					ca( 51) <= SEED( 43) xor SEED(185) xor SEED(186) xor SEED(190) xor dq( 51);
					ca( 52) <= SEED( 44) xor SEED(186) xor SEED(187) xor SEED(191) xor dq( 52);
					ca( 53) <= SEED( 45) xor SEED(187) xor SEED(188) xor dq( 53);
					ca( 54) <= SEED( 46) xor SEED(184) xor SEED(186) xor SEED(191) xor dq( 54);
					ca( 55) <= SEED( 47) xor SEED(185) xor SEED(187) xor dq( 55);
					ca( 56) <= SEED( 48) xor SEED(184) xor SEED(189) xor SEED(191) xor dq( 56);
					ca( 57) <= SEED( 49) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 57);
					ca( 58) <= SEED( 50) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 58);
					ca( 59) <= SEED( 51) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq( 59);
					ca( 60) <= SEED( 52) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq( 60);
					ca( 61) <= SEED( 53) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 61);
					ca( 62) <= SEED( 54) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 62);
					ca( 63) <= SEED( 55) xor SEED(190) xor SEED(191) xor dq( 63);
					ca( 64) <= SEED( 56) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor dq( 64);
					ca( 65) <= SEED( 57) xor SEED(185) xor SEED(187) xor SEED(189) xor SEED(190) xor dq( 65);
					ca( 66) <= SEED( 58) xor SEED(186) xor SEED(188) xor SEED(190) xor SEED(191) xor dq( 66);
					ca( 67) <= SEED( 59) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(188) xor dq( 67);
					ca( 68) <= SEED( 60) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(189) xor dq( 68);
					ca( 69) <= SEED( 61) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 69);
					ca( 70) <= SEED( 62) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 70);
					ca( 71) <= SEED( 63) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(190) xor dq( 71);
					ca( 72) <= SEED( 64) xor SEED(185) xor SEED(187) xor SEED(190) xor SEED(191) xor dq( 72);
					ca( 73) <= SEED( 65) xor SEED(186) xor SEED(188) xor SEED(191) xor dq( 73);
					ca( 74) <= SEED( 66) xor SEED(187) xor SEED(189) xor dq( 74);
					ca( 75) <= SEED( 67) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 75);
					ca( 76) <= SEED( 68) xor SEED(185) xor SEED(187) xor SEED(190) xor SEED(191) xor dq( 76);
					ca( 77) <= SEED( 69) xor SEED(186) xor SEED(188) xor SEED(191) xor dq( 77);
					ca( 78) <= SEED( 70) xor SEED(187) xor SEED(189) xor dq( 78);
					ca( 79) <= SEED( 71) xor SEED(188) xor SEED(190) xor dq( 79);
					ca( 80) <= SEED( 72) xor SEED(184) xor SEED(186) xor SEED(188) xor dq( 80);
					ca( 81) <= SEED( 73) xor SEED(185) xor SEED(187) xor SEED(189) xor dq( 81);
					ca( 82) <= SEED( 74) xor SEED(184) xor SEED(189) xor SEED(190) xor SEED(191) xor dq( 82);
					ca( 83) <= SEED( 75) xor SEED(185) xor SEED(190) xor SEED(191) xor dq( 83);
					ca( 84) <= SEED( 76) xor SEED(184) xor SEED(188) xor SEED(189) xor dq( 84);
					ca( 85) <= SEED( 77) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(190) xor SEED(191) xor dq( 85);
					ca( 86) <= SEED( 78) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(191) xor dq( 86);
					ca( 87) <= SEED( 79) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor dq( 87);
					ca( 88) <= SEED( 80) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq( 88);
					ca( 89) <= SEED( 81) xor SEED(188) xor SEED(189) xor SEED(190) xor dq( 89);
					ca( 90) <= SEED( 82) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(190) xor dq( 90);
					ca( 91) <= SEED( 83) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor dq( 91);
					ca( 92) <= SEED( 84) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(191) xor dq( 92);
					ca( 93) <= SEED( 85) xor SEED(185) xor SEED(186) xor SEED(188) xor dq( 93);
					ca( 94) <= SEED( 86) xor SEED(184) xor SEED(187) xor SEED(188) xor SEED(191) xor dq( 94);
					ca( 95) <= SEED( 87) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(191) xor dq( 95);
					ca( 96) <= SEED( 88) xor SEED(185) xor SEED(186) xor SEED(187) xor dq( 96);
					ca( 97) <= SEED( 89) xor SEED(186) xor SEED(187) xor SEED(188) xor dq( 97);
					ca( 98) <= SEED( 90) xor SEED(187) xor SEED(188) xor SEED(189) xor dq( 98);
					ca( 99) <= SEED( 91) xor SEED(184) xor SEED(186) xor SEED(190) xor SEED(191) xor dq( 99);
					ca(100) <= SEED( 92) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor dq(100);
					ca(101) <= SEED( 93) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(101);
					ca(102) <= SEED( 94) xor SEED(184) xor SEED(187) xor SEED(190) xor dq(102);
					ca(103) <= SEED( 95) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(189) xor dq(103);
					ca(104) <= SEED( 96) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(190) xor dq(104);
					ca(105) <= SEED( 97) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(191) xor dq(105);
					ca(106) <= SEED( 98) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(191) xor dq(106);
					ca(107) <= SEED( 99) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(191) xor dq(107);
					ca(108) <= SEED(100) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor dq(108);
					ca(109) <= SEED(101) xor SEED(184) xor SEED(187) xor dq(109);
					ca(110) <= SEED(102) xor SEED(185) xor SEED(188) xor dq(110);
					ca(111) <= SEED(103) xor SEED(186) xor SEED(189) xor dq(111);
					ca(112) <= SEED(104) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(112);
					ca(113) <= SEED(105) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(190) xor dq(113);
					ca(114) <= SEED(106) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(189) xor dq(114);
					ca(115) <= SEED(107) xor SEED(184) xor SEED(185) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(115);
					ca(116) <= SEED(108) xor SEED(185) xor SEED(186) xor SEED(190) xor SEED(191) xor dq(116);
					ca(117) <= SEED(109) xor SEED(186) xor SEED(187) xor SEED(191) xor dq(117);
					ca(118) <= SEED(110) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(191) xor dq(118);
					ca(119) <= SEED(111) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(119);
					ca(120) <= SEED(112) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq(120);
					ca(121) <= SEED(113) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(121);
					ca(122) <= SEED(114) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(122);
					ca(123) <= SEED(115) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(123);
					ca(124) <= SEED(116) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(190) xor dq(124);
					ca(125) <= SEED(117) xor SEED(185) xor SEED(187) xor SEED(189) xor SEED(191) xor dq(125);
					ca(126) <= SEED(118) xor SEED(184) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(126);
					ca(127) <= SEED(119) xor SEED(185) xor SEED(190) xor SEED(191) xor dq(127);
					ca(128) <= SEED(120) xor SEED(186) xor SEED(191) xor dq(128);
					ca(129) <= SEED(121) xor SEED(187) xor dq(129);
					ca(130) <= SEED(122) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(191) xor dq(130);
					ca(131) <= SEED(123) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(131);
					ca(132) <= SEED(124) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(190) xor dq(132);
					ca(133) <= SEED(125) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(191) xor dq(133);
					ca(134) <= SEED(126) xor SEED(186) xor SEED(187) xor SEED(189) xor dq(134);
					ca(135) <= SEED(127) xor SEED(187) xor SEED(188) xor SEED(190) xor dq(135);
					ca(136) <= SEED(128) xor SEED(184) xor SEED(186) xor dq(136);
					ca(137) <= SEED(129) xor SEED(185) xor SEED(187) xor dq(137);
					ca(138) <= SEED(130) xor SEED(186) xor SEED(188) xor dq(138);
					ca(139) <= SEED(131) xor SEED(187) xor SEED(189) xor dq(139);
					ca(140) <= SEED(132) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(140);
					ca(141) <= SEED(133) xor SEED(185) xor SEED(187) xor SEED(190) xor SEED(191) xor dq(141);
					ca(142) <= SEED(134) xor SEED(184) xor SEED(189) xor dq(142);
					ca(143) <= SEED(135) xor SEED(185) xor SEED(190) xor dq(143);
					ca(144) <= SEED(136) xor SEED(186) xor SEED(191) xor dq(144);
					ca(145) <= SEED(137) xor SEED(187) xor dq(145);
					ca(146) <= SEED(138) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(191) xor dq(146);
					ca(147) <= SEED(139) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(147);
					ca(148) <= SEED(140) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(190) xor dq(148);
					ca(149) <= SEED(141) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(191) xor dq(149);
					ca(150) <= SEED(142) xor SEED(184) xor SEED(187) xor SEED(188) xor SEED(191) xor dq(150);
					ca(151) <= SEED(143) xor SEED(185) xor SEED(188) xor SEED(189) xor dq(151);
					ca(152) <= SEED(144) xor SEED(186) xor SEED(189) xor SEED(190) xor dq(152);
					ca(153) <= SEED(145) xor SEED(187) xor SEED(190) xor SEED(191) xor dq(153);
					ca(154) <= SEED(146) xor SEED(184) xor SEED(186) xor SEED(189) xor dq(154);
					ca(155) <= SEED(147) xor SEED(185) xor SEED(187) xor SEED(190) xor dq(155);
					ca(156) <= SEED(148) xor SEED(186) xor SEED(188) xor SEED(191) xor dq(156);
					ca(157) <= SEED(149) xor SEED(187) xor SEED(189) xor dq(157);
					ca(158) <= SEED(150) xor SEED(188) xor SEED(190) xor dq(158);
					ca(159) <= SEED(151) xor SEED(184) xor SEED(186) xor SEED(188) xor dq(159);
					ca(160) <= SEED(152) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(191) xor dq(160);
					ca(161) <= SEED(153) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(191) xor dq(161);
					ca(162) <= SEED(154) xor SEED(185) xor SEED(186) xor SEED(188) xor dq(162);
					ca(163) <= SEED(155) xor SEED(186) xor SEED(187) xor SEED(189) xor dq(163);
					ca(164) <= SEED(156) xor SEED(187) xor SEED(188) xor SEED(190) xor dq(164);
					ca(165) <= SEED(157) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(165);
					ca(166) <= SEED(158) xor SEED(189) xor SEED(190) xor dq(166);
					ca(167) <= SEED(159) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(167);
					ca(168) <= SEED(160) xor SEED(185) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(168);
					ca(169) <= SEED(161) xor SEED(184) xor SEED(189) xor SEED(190) xor dq(169);
					ca(170) <= SEED(162) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(170);
					ca(171) <= SEED(163) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(190) xor dq(171);
					ca(172) <= SEED(164) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(172);
					ca(173) <= SEED(165) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor dq(173);
					ca(174) <= SEED(166) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq(174);
					ca(175) <= SEED(167) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(175);
					ca(176) <= SEED(168) xor SEED(189) xor SEED(190) xor dq(176);
					ca(177) <= SEED(169) xor SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(177);
					ca(178) <= SEED(170) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(190) xor dq(178);
					ca(179) <= SEED(171) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(179);
					ca(180) <= SEED(172) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(180);
					ca(181) <= SEED(173) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(190) xor dq(181);
					ca(182) <= SEED(174) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(191) xor dq(182);
					ca(183) <= SEED(175) xor SEED(186) xor SEED(188) xor SEED(189) xor dq(183);
					ca(184) <= SEED(176) xor SEED(187) xor SEED(189) xor SEED(190) xor dq(184);
					ca(185) <= SEED(177) xor SEED(184) xor SEED(186) xor SEED(189) xor SEED(190) xor dq(185);
					ca(186) <= SEED(178) xor SEED(184) xor SEED(185) xor SEED(186) xor SEED(187) xor SEED(188) xor SEED(189) xor SEED(190) xor dq(186);
					ca(187) <= SEED(179) xor SEED(184) xor SEED(185) xor SEED(187) xor SEED(190) xor dq(187);
					ca(188) <= SEED(180) xor SEED(185) xor SEED(186) xor SEED(188) xor SEED(191) xor dq(188);
					ca(189) <= SEED(181) xor SEED(186) xor SEED(187) xor SEED(189) xor dq(189);
					ca(190) <= SEED(182) xor SEED(184) xor SEED(186) xor SEED(187) xor SEED(189) xor SEED(190) xor SEED(191) xor dq(190);
					ca(191) <= SEED(183) xor SEED(185) xor SEED(187) xor SEED(188) xor SEED(190) xor SEED(191) xor dq(191);


					oa(  7) <= SEED(191) xor dq(  0);
					oa(  6) <= SEED(190) xor dq(  1);
					oa(  5) <= SEED(189) xor SEED(191) xor dq(  2);
					oa(  4) <= SEED(188) xor SEED(190) xor dq(  3);
					oa(  3) <= SEED(187) xor SEED(189) xor SEED(191) xor dq(  4);
					oa(  2) <= SEED(186) xor SEED(188) xor SEED(190) xor SEED(191) xor dq(  5);
					oa(  1) <= SEED(185) xor SEED(187) xor SEED(189) xor SEED(190) xor dq(  6);
					oa(  0) <= SEED(184) xor SEED(186) xor SEED(188) xor SEED(189) xor SEED(191) xor dq(  7);
				else
					ca(  0) <= ca(184) xor ca(186) xor ca(188) xor ca(189) xor ca(191) xor dq(  0);
					ca(  1) <= ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq(  1);
					ca(  2) <= ca(184) xor ca(185) xor ca(187) xor dq(  2);
					ca(  3) <= ca(185) xor ca(186) xor ca(188) xor dq(  3);
					ca(  4) <= ca(186) xor ca(187) xor ca(189) xor dq(  4);
					ca(  5) <= ca(184) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq(  5);
					ca(  6) <= ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor dq(  6);
					ca(  7) <= ca(184) xor ca(185) xor ca(187) xor ca(189) xor ca(190) xor dq(  7);
					ca(  8) <= ca(  0) xor ca(184) xor ca(185) xor ca(189) xor ca(190) xor dq(  8);
					ca(  9) <= ca(  1) xor ca(185) xor ca(186) xor ca(190) xor ca(191) xor dq(  9);
					ca( 10) <= ca(  2) xor ca(184) xor ca(187) xor ca(188) xor ca(189) xor dq( 10);
					ca( 11) <= ca(  3) xor ca(185) xor ca(188) xor ca(189) xor ca(190) xor dq( 11);
					ca( 12) <= ca(  4) xor ca(184) xor ca(188) xor ca(190) xor dq( 12);
					ca( 13) <= ca(  5) xor ca(185) xor ca(189) xor ca(191) xor dq( 13);
					ca( 14) <= ca(  6) xor ca(184) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 14);
					ca( 15) <= ca(  7) xor ca(185) xor ca(189) xor ca(190) xor ca(191) xor dq( 15);
					ca( 16) <= ca(  8) xor ca(186) xor ca(190) xor ca(191) xor dq( 16);
					ca( 17) <= ca(  9) xor ca(184) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor dq( 17);
					ca( 18) <= ca( 10) xor ca(185) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq( 18);
					ca( 19) <= ca( 11) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 19);
					ca( 20) <= ca( 12) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq( 20);
					ca( 21) <= ca( 13) xor ca(188) xor ca(190) xor ca(191) xor dq( 21);
					ca( 22) <= ca( 14) xor ca(189) xor ca(191) xor dq( 22);
					ca( 23) <= ca( 15) xor ca(190) xor dq( 23);
					ca( 24) <= ca( 16) xor ca(191) xor dq( 24);
					ca( 25) <= ca( 17) xor ca(184) xor ca(186) xor ca(188) xor ca(189) xor ca(191) xor dq( 25);
					ca( 26) <= ca( 18) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq( 26);
					ca( 27) <= ca( 19) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq( 27);
					ca( 28) <= ca( 20) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq( 28);
					ca( 29) <= ca( 21) xor ca(184) xor ca(186) xor ca(187) xor ca(190) xor dq( 29);
					ca( 30) <= ca( 22) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor dq( 30);
					ca( 31) <= ca( 23) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor dq( 31);
					ca( 32) <= ca( 24) xor ca(184) xor ca(187) xor dq( 32);
					ca( 33) <= ca( 25) xor ca(184) xor ca(185) xor ca(186) xor ca(189) xor ca(191) xor dq( 33);
					ca( 34) <= ca( 26) xor ca(184) xor ca(185) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 34);
					ca( 35) <= ca( 27) xor ca(185) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 35);
					ca( 36) <= ca( 28) xor ca(184) xor ca(187) xor ca(188) xor ca(190) xor dq( 36);
					ca( 37) <= ca( 29) xor ca(184) xor ca(185) xor ca(186) xor dq( 37);
					ca( 38) <= ca( 30) xor ca(184) xor ca(185) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq( 38);
					ca( 39) <= ca( 31) xor ca(184) xor ca(185) xor ca(190) xor ca(191) xor dq( 39);
					ca( 40) <= ca( 32) xor ca(184) xor ca(185) xor ca(188) xor ca(189) xor dq( 40);
					ca( 41) <= ca( 33) xor ca(185) xor ca(186) xor ca(189) xor ca(190) xor dq( 41);
					ca( 42) <= ca( 34) xor ca(184) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq( 42);
					ca( 43) <= ca( 35) xor ca(185) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 43);
					ca( 44) <= ca( 36) xor ca(186) xor ca(189) xor ca(190) xor ca(191) xor dq( 44);
					ca( 45) <= ca( 37) xor ca(187) xor ca(190) xor ca(191) xor dq( 45);
					ca( 46) <= ca( 38) xor ca(188) xor ca(191) xor dq( 46);
					ca( 47) <= ca( 39) xor ca(184) xor ca(186) xor ca(188) xor ca(191) xor dq( 47);
					ca( 48) <= ca( 40) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(191) xor dq( 48);
					ca( 49) <= ca( 41) xor ca(184) xor ca(185) xor ca(187) xor ca(191) xor dq( 49);
					ca( 50) <= ca( 42) xor ca(184) xor ca(185) xor ca(189) xor ca(191) xor dq( 50);
					ca( 51) <= ca( 43) xor ca(185) xor ca(186) xor ca(190) xor dq( 51);
					ca( 52) <= ca( 44) xor ca(186) xor ca(187) xor ca(191) xor dq( 52);
					ca( 53) <= ca( 45) xor ca(187) xor ca(188) xor dq( 53);
					ca( 54) <= ca( 46) xor ca(184) xor ca(186) xor ca(191) xor dq( 54);
					ca( 55) <= ca( 47) xor ca(185) xor ca(187) xor dq( 55);
					ca( 56) <= ca( 48) xor ca(184) xor ca(189) xor ca(191) xor dq( 56);
					ca( 57) <= ca( 49) xor ca(184) xor ca(185) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq( 57);
					ca( 58) <= ca( 50) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq( 58);
					ca( 59) <= ca( 51) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq( 59);
					ca( 60) <= ca( 52) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq( 60);
					ca( 61) <= ca( 53) xor ca(188) xor ca(189) xor ca(190) xor dq( 61);
					ca( 62) <= ca( 54) xor ca(189) xor ca(190) xor ca(191) xor dq( 62);
					ca( 63) <= ca( 55) xor ca(190) xor ca(191) xor dq( 63);
					ca( 64) <= ca( 56) xor ca(184) xor ca(186) xor ca(188) xor ca(189) xor dq( 64);
					ca( 65) <= ca( 57) xor ca(185) xor ca(187) xor ca(189) xor ca(190) xor dq( 65);
					ca( 66) <= ca( 58) xor ca(186) xor ca(188) xor ca(190) xor ca(191) xor dq( 66);
					ca( 67) <= ca( 59) xor ca(184) xor ca(186) xor ca(187) xor ca(188) xor dq( 67);
					ca( 68) <= ca( 60) xor ca(185) xor ca(187) xor ca(188) xor ca(189) xor dq( 68);
					ca( 69) <= ca( 61) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor dq( 69);
					ca( 70) <= ca( 62) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq( 70);
					ca( 71) <= ca( 63) xor ca(184) xor ca(186) xor ca(189) xor ca(190) xor dq( 71);
					ca( 72) <= ca( 64) xor ca(185) xor ca(187) xor ca(190) xor ca(191) xor dq( 72);
					ca( 73) <= ca( 65) xor ca(186) xor ca(188) xor ca(191) xor dq( 73);
					ca( 74) <= ca( 66) xor ca(187) xor ca(189) xor dq( 74);
					ca( 75) <= ca( 67) xor ca(184) xor ca(186) xor ca(189) xor ca(190) xor ca(191) xor dq( 75);
					ca( 76) <= ca( 68) xor ca(185) xor ca(187) xor ca(190) xor ca(191) xor dq( 76);
					ca( 77) <= ca( 69) xor ca(186) xor ca(188) xor ca(191) xor dq( 77);
					ca( 78) <= ca( 70) xor ca(187) xor ca(189) xor dq( 78);
					ca( 79) <= ca( 71) xor ca(188) xor ca(190) xor dq( 79);
					ca( 80) <= ca( 72) xor ca(184) xor ca(186) xor ca(188) xor dq( 80);
					ca( 81) <= ca( 73) xor ca(185) xor ca(187) xor ca(189) xor dq( 81);
					ca( 82) <= ca( 74) xor ca(184) xor ca(189) xor ca(190) xor ca(191) xor dq( 82);
					ca( 83) <= ca( 75) xor ca(185) xor ca(190) xor ca(191) xor dq( 83);
					ca( 84) <= ca( 76) xor ca(184) xor ca(188) xor ca(189) xor dq( 84);
					ca( 85) <= ca( 77) xor ca(184) xor ca(185) xor ca(186) xor ca(188) xor ca(190) xor ca(191) xor dq( 85);
					ca( 86) <= ca( 78) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor ca(191) xor dq( 86);
					ca( 87) <= ca( 79) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor dq( 87);
					ca( 88) <= ca( 80) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq( 88);
					ca( 89) <= ca( 81) xor ca(188) xor ca(189) xor ca(190) xor dq( 89);
					ca( 90) <= ca( 82) xor ca(184) xor ca(186) xor ca(188) xor ca(190) xor dq( 90);
					ca( 91) <= ca( 83) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor dq( 91);
					ca( 92) <= ca( 84) xor ca(184) xor ca(185) xor ca(187) xor ca(191) xor dq( 92);
					ca( 93) <= ca( 85) xor ca(185) xor ca(186) xor ca(188) xor dq( 93);
					ca( 94) <= ca( 86) xor ca(184) xor ca(187) xor ca(188) xor ca(191) xor dq( 94);
					ca( 95) <= ca( 87) xor ca(184) xor ca(185) xor ca(186) xor ca(191) xor dq( 95);
					ca( 96) <= ca( 88) xor ca(185) xor ca(186) xor ca(187) xor dq( 96);
					ca( 97) <= ca( 89) xor ca(186) xor ca(187) xor ca(188) xor dq( 97);
					ca( 98) <= ca( 90) xor ca(187) xor ca(188) xor ca(189) xor dq( 98);
					ca( 99) <= ca( 91) xor ca(184) xor ca(186) xor ca(190) xor ca(191) xor dq( 99);
					ca(100) <= ca( 92) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor dq(100);
					ca(101) <= ca( 93) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq(101);
					ca(102) <= ca( 94) xor ca(184) xor ca(187) xor ca(190) xor dq(102);
					ca(103) <= ca( 95) xor ca(184) xor ca(185) xor ca(186) xor ca(189) xor dq(103);
					ca(104) <= ca( 96) xor ca(185) xor ca(186) xor ca(187) xor ca(190) xor dq(104);
					ca(105) <= ca( 97) xor ca(186) xor ca(187) xor ca(188) xor ca(191) xor dq(105);
					ca(106) <= ca( 98) xor ca(184) xor ca(186) xor ca(187) xor ca(191) xor dq(106);
					ca(107) <= ca( 99) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor ca(191) xor dq(107);
					ca(108) <= ca(100) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor dq(108);
					ca(109) <= ca(101) xor ca(184) xor ca(187) xor dq(109);
					ca(110) <= ca(102) xor ca(185) xor ca(188) xor dq(110);
					ca(111) <= ca(103) xor ca(186) xor ca(189) xor dq(111);
					ca(112) <= ca(104) xor ca(184) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq(112);
					ca(113) <= ca(105) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(190) xor dq(113);
					ca(114) <= ca(106) xor ca(184) xor ca(185) xor ca(187) xor ca(189) xor dq(114);
					ca(115) <= ca(107) xor ca(184) xor ca(185) xor ca(189) xor ca(190) xor ca(191) xor dq(115);
					ca(116) <= ca(108) xor ca(185) xor ca(186) xor ca(190) xor ca(191) xor dq(116);
					ca(117) <= ca(109) xor ca(186) xor ca(187) xor ca(191) xor dq(117);
					ca(118) <= ca(110) xor ca(184) xor ca(186) xor ca(187) xor ca(189) xor ca(191) xor dq(118);
					ca(119) <= ca(111) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq(119);
					ca(120) <= ca(112) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq(120);
					ca(121) <= ca(113) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq(121);
					ca(122) <= ca(114) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq(122);
					ca(123) <= ca(115) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq(123);
					ca(124) <= ca(116) xor ca(184) xor ca(186) xor ca(188) xor ca(190) xor dq(124);
					ca(125) <= ca(117) xor ca(185) xor ca(187) xor ca(189) xor ca(191) xor dq(125);
					ca(126) <= ca(118) xor ca(184) xor ca(189) xor ca(190) xor ca(191) xor dq(126);
					ca(127) <= ca(119) xor ca(185) xor ca(190) xor ca(191) xor dq(127);
					ca(128) <= ca(120) xor ca(186) xor ca(191) xor dq(128);
					ca(129) <= ca(121) xor ca(187) xor dq(129);
					ca(130) <= ca(122) xor ca(184) xor ca(186) xor ca(189) xor ca(191) xor dq(130);
					ca(131) <= ca(123) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq(131);
					ca(132) <= ca(124) xor ca(184) xor ca(185) xor ca(187) xor ca(190) xor dq(132);
					ca(133) <= ca(125) xor ca(185) xor ca(186) xor ca(188) xor ca(191) xor dq(133);
					ca(134) <= ca(126) xor ca(186) xor ca(187) xor ca(189) xor dq(134);
					ca(135) <= ca(127) xor ca(187) xor ca(188) xor ca(190) xor dq(135);
					ca(136) <= ca(128) xor ca(184) xor ca(186) xor dq(136);
					ca(137) <= ca(129) xor ca(185) xor ca(187) xor dq(137);
					ca(138) <= ca(130) xor ca(186) xor ca(188) xor dq(138);
					ca(139) <= ca(131) xor ca(187) xor ca(189) xor dq(139);
					ca(140) <= ca(132) xor ca(184) xor ca(186) xor ca(189) xor ca(190) xor ca(191) xor dq(140);
					ca(141) <= ca(133) xor ca(185) xor ca(187) xor ca(190) xor ca(191) xor dq(141);
					ca(142) <= ca(134) xor ca(184) xor ca(189) xor dq(142);
					ca(143) <= ca(135) xor ca(185) xor ca(190) xor dq(143);
					ca(144) <= ca(136) xor ca(186) xor ca(191) xor dq(144);
					ca(145) <= ca(137) xor ca(187) xor dq(145);
					ca(146) <= ca(138) xor ca(184) xor ca(186) xor ca(189) xor ca(191) xor dq(146);
					ca(147) <= ca(139) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor ca(191) xor dq(147);
					ca(148) <= ca(140) xor ca(184) xor ca(185) xor ca(187) xor ca(190) xor dq(148);
					ca(149) <= ca(141) xor ca(185) xor ca(186) xor ca(188) xor ca(191) xor dq(149);
					ca(150) <= ca(142) xor ca(184) xor ca(187) xor ca(188) xor ca(191) xor dq(150);
					ca(151) <= ca(143) xor ca(185) xor ca(188) xor ca(189) xor dq(151);
					ca(152) <= ca(144) xor ca(186) xor ca(189) xor ca(190) xor dq(152);
					ca(153) <= ca(145) xor ca(187) xor ca(190) xor ca(191) xor dq(153);
					ca(154) <= ca(146) xor ca(184) xor ca(186) xor ca(189) xor dq(154);
					ca(155) <= ca(147) xor ca(185) xor ca(187) xor ca(190) xor dq(155);
					ca(156) <= ca(148) xor ca(186) xor ca(188) xor ca(191) xor dq(156);
					ca(157) <= ca(149) xor ca(187) xor ca(189) xor dq(157);
					ca(158) <= ca(150) xor ca(188) xor ca(190) xor dq(158);
					ca(159) <= ca(151) xor ca(184) xor ca(186) xor ca(188) xor dq(159);
					ca(160) <= ca(152) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(191) xor dq(160);
					ca(161) <= ca(153) xor ca(184) xor ca(185) xor ca(187) xor ca(191) xor dq(161);
					ca(162) <= ca(154) xor ca(185) xor ca(186) xor ca(188) xor dq(162);
					ca(163) <= ca(155) xor ca(186) xor ca(187) xor ca(189) xor dq(163);
					ca(164) <= ca(156) xor ca(187) xor ca(188) xor ca(190) xor dq(164);
					ca(165) <= ca(157) xor ca(188) xor ca(189) xor ca(191) xor dq(165);
					ca(166) <= ca(158) xor ca(189) xor ca(190) xor dq(166);
					ca(167) <= ca(159) xor ca(184) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor dq(167);
					ca(168) <= ca(160) xor ca(185) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq(168);
					ca(169) <= ca(161) xor ca(184) xor ca(189) xor ca(190) xor dq(169);
					ca(170) <= ca(162) xor ca(184) xor ca(185) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor dq(170);
					ca(171) <= ca(163) xor ca(184) xor ca(185) xor ca(187) xor ca(188) xor ca(190) xor dq(171);
					ca(172) <= ca(164) xor ca(185) xor ca(186) xor ca(188) xor ca(189) xor ca(191) xor dq(172);
					ca(173) <= ca(165) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor dq(173);
					ca(174) <= ca(166) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq(174);
					ca(175) <= ca(167) xor ca(188) xor ca(189) xor ca(191) xor dq(175);
					ca(176) <= ca(168) xor ca(189) xor ca(190) xor dq(176);
					ca(177) <= ca(169) xor ca(184) xor ca(186) xor ca(188) xor ca(189) xor ca(190) xor dq(177);
					ca(178) <= ca(170) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(190) xor dq(178);
					ca(179) <= ca(171) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(191) xor dq(179);
					ca(180) <= ca(172) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq(180);
					ca(181) <= ca(173) xor ca(184) xor ca(186) xor ca(187) xor ca(190) xor dq(181);
					ca(182) <= ca(174) xor ca(185) xor ca(187) xor ca(188) xor ca(191) xor dq(182);
					ca(183) <= ca(175) xor ca(186) xor ca(188) xor ca(189) xor dq(183);
					ca(184) <= ca(176) xor ca(187) xor ca(189) xor ca(190) xor dq(184);
					ca(185) <= ca(177) xor ca(184) xor ca(186) xor ca(189) xor ca(190) xor dq(185);
					ca(186) <= ca(178) xor ca(184) xor ca(185) xor ca(186) xor ca(187) xor ca(188) xor ca(189) xor ca(190) xor dq(186);
					ca(187) <= ca(179) xor ca(184) xor ca(185) xor ca(187) xor ca(190) xor dq(187);
					ca(188) <= ca(180) xor ca(185) xor ca(186) xor ca(188) xor ca(191) xor dq(188);
					ca(189) <= ca(181) xor ca(186) xor ca(187) xor ca(189) xor dq(189);
					ca(190) <= ca(182) xor ca(184) xor ca(186) xor ca(187) xor ca(189) xor ca(190) xor ca(191) xor dq(190);
					ca(191) <= ca(183) xor ca(185) xor ca(187) xor ca(188) xor ca(190) xor ca(191) xor dq(191);


					oa(  7) <= ca(191) xor dq(  0);
					oa(  6) <= ca(190) xor dq(  1);
					oa(  5) <= ca(189) xor ca(191) xor dq(  2);
					oa(  4) <= ca(188) xor ca(190) xor dq(  3);
					oa(  3) <= ca(187) xor ca(189) xor ca(191) xor dq(  4);
					oa(  2) <= ca(186) xor ca(188) xor ca(190) xor ca(191) xor dq(  5);
					oa(  1) <= ca(185) xor ca(187) xor ca(189) xor ca(190) xor dq(  6);
					oa(  0) <= ca(184) xor ca(186) xor ca(188) xor ca(189) xor ca(191) xor dq(  7);
				end if;
			end if;
		end if;
	end process;
	c <= ca;
	o <= oa;
end a1;
