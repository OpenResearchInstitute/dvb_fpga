--
-- DVB IP
--
-- Copyright 2020 by Suoto <andre820@gmail.com>
--
-- This file is part of the DVB IP.
--
-- DVB IP is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- DVB IP is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with DVB IP.  If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library fpga_cores;
use fpga_cores.common_pkg.all;

use work.dvb_utils_pkg.all;

-- Summary of statistics

--    table                               depth    width (bits)    width (entries)    total (bytes)    18k BRAMs    36k BRAMs
----  --------------------------------  -------  --------------  -----------------  ---------------  -----------  -----------
--    ldpc_table_FECFRAME_NORMAL_C1_2        90             115                  9             1294            7            4
--    ldpc_table_FECFRAME_NORMAL_C1_3        60             196                 13             1470           11            6
--    ldpc_table_FECFRAME_NORMAL_C1_4        45             196                 13             1103           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_3       120             189                 14             2835           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_5        72             196                 13             1764           11            6
--    ldpc_table_FECFRAME_NORMAL_C3_4       135             164                 13             2768           10            5
--    ldpc_table_FECFRAME_NORMAL_C3_5       108             184                 13             2484           11            6
--    ldpc_table_FECFRAME_NORMAL_C4_5       144             150                 12             2700            9            5
--    ldpc_table_FECFRAME_NORMAL_C5_6       150             177                 14             3319           10            5
--    ldpc_table_FECFRAME_NORMAL_C8_9       160              46                  5              920            3            2
--    ldpc_table_FECFRAME_NORMAL_C9_10      162              46                  5              932            3            2
--    ldpc_table_FECFRAME_SHORT_C1_2         20             100                  9              250            6            3
--    ldpc_table_FECFRAME_SHORT_C1_3         15             170                 13              319           10            5
--    ldpc_table_FECFRAME_SHORT_C1_4          9             171                 13              193           10            5
--    ldpc_table_FECFRAME_SHORT_C2_3         30             156                 14              585            9            5
--    ldpc_table_FECFRAME_SHORT_C2_5         18             168                 13              378           10            5
--    ldpc_table_FECFRAME_SHORT_C3_4         33             133                 13              549            8            4
--    ldpc_table_FECFRAME_SHORT_C3_5         27             160                 13              540            9            5
--    ldpc_table_FECFRAME_SHORT_C4_5         35              30                  4              132            2            1
--    ldpc_table_FECFRAME_SHORT_C5_6         37             139                 14              643            8            4
--    ldpc_table_FECFRAME_SHORT_C8_9         40              37                  5              185            3            2

package ldpc_tables_pkg is


  -- LDPC_TABLE_FECFRAME_<frame_length>_<code_rate>_COLUMN_WIDTHS constants have the bit
  -- width of each row

  -- LDPC_TABLE_FECFRAME_<frame_length>_<code_rate> is the actual LDPC where the number of
  -- columns is normalized to the row with most columns and the first column of each row
  -- contains the number of valid elements within the row. Elements outisde the valid range
  -- are represented as -1


  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_2.csv, table is 90x115 (1293.75 bytes)
  -- Resource estimation: 7 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 7, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2 : integer_2d_array_t(0 to 89)(0 to 8) := (
    0 => integer_vector_t'(0 => 8, 1 => 54, 2 => 9318, 3 => 14392, 4 => 27561, 5 => 26909, 6 => 10219, 7 => 2534, 8 => 8597),
    1 => integer_vector_t'(0 => 8, 1 => 55, 2 => 7263, 3 => 4635, 4 => 2530, 5 => 28130, 6 => 3033, 7 => 23830, 8 => 3651),
    2 => integer_vector_t'(0 => 8, 1 => 56, 2 => 24731, 3 => 23583, 4 => 26036, 5 => 17299, 6 => 5750, 7 => 792, 8 => 9169),
    3 => integer_vector_t'(0 => 8, 1 => 57, 2 => 5811, 3 => 26154, 4 => 18653, 5 => 11551, 6 => 15447, 7 => 13685, 8 => 16264),
    4 => integer_vector_t'(0 => 8, 1 => 58, 2 => 12610, 3 => 11347, 4 => 28768, 5 => 2792, 6 => 3174, 7 => 29371, 8 => 12997),
    5 => integer_vector_t'(0 => 8, 1 => 59, 2 => 16789, 3 => 16018, 4 => 21449, 5 => 6165, 6 => 21202, 7 => 15850, 8 => 3186),
    6 => integer_vector_t'(0 => 8, 1 => 60, 2 => 31016, 3 => 21449, 4 => 17618, 5 => 6213, 6 => 12166, 7 => 8334, 8 => 18212),
    7 => integer_vector_t'(0 => 8, 1 => 61, 2 => 22836, 3 => 14213, 4 => 11327, 5 => 5896, 6 => 718, 7 => 11727, 8 => 9308),
    8 => integer_vector_t'(0 => 8, 1 => 62, 2 => 2091, 3 => 24941, 4 => 29966, 5 => 23634, 6 => 9013, 7 => 15587, 8 => 5444),
    9 => integer_vector_t'(0 => 8, 1 => 63, 2 => 22207, 3 => 3983, 4 => 16904, 5 => 28534, 6 => 21415, 7 => 27524, 8 => 25912),
    10 => integer_vector_t'(0 => 8, 1 => 64, 2 => 25687, 3 => 4501, 4 => 22193, 5 => 14665, 6 => 14798, 7 => 16158, 8 => 5491),
    11 => integer_vector_t'(0 => 8, 1 => 65, 2 => 4520, 3 => 17094, 4 => 23397, 5 => 4264, 6 => 22370, 7 => 16941, 8 => 21526),
    12 => integer_vector_t'(0 => 8, 1 => 66, 2 => 10490, 3 => 6182, 4 => 32370, 5 => 9597, 6 => 30841, 7 => 25954, 8 => 2762),
    13 => integer_vector_t'(0 => 8, 1 => 67, 2 => 22120, 3 => 22865, 4 => 29870, 5 => 15147, 6 => 13668, 7 => 14955, 8 => 19235),
    14 => integer_vector_t'(0 => 8, 1 => 68, 2 => 6689, 3 => 18408, 4 => 18346, 5 => 9918, 6 => 25746, 7 => 5443, 8 => 20645),
    15 => integer_vector_t'(0 => 8, 1 => 69, 2 => 29982, 3 => 12529, 4 => 13858, 5 => 4746, 6 => 30370, 7 => 10023, 8 => 24828),
    16 => integer_vector_t'(0 => 8, 1 => 70, 2 => 1262, 3 => 28032, 4 => 29888, 5 => 13063, 6 => 24033, 7 => 21951, 8 => 7863),
    17 => integer_vector_t'(0 => 8, 1 => 71, 2 => 6594, 3 => 29642, 4 => 31451, 5 => 14831, 6 => 9509, 7 => 9335, 8 => 31552),
    18 => integer_vector_t'(0 => 8, 1 => 72, 2 => 1358, 3 => 6454, 4 => 16633, 5 => 20354, 6 => 24598, 7 => 624, 8 => 5265),
    19 => integer_vector_t'(0 => 8, 1 => 73, 2 => 19529, 3 => 295, 4 => 18011, 5 => 3080, 6 => 13364, 7 => 8032, 8 => 15323),
    20 => integer_vector_t'(0 => 8, 1 => 74, 2 => 11981, 3 => 1510, 4 => 7960, 5 => 21462, 6 => 9129, 7 => 11370, 8 => 25741),
    21 => integer_vector_t'(0 => 8, 1 => 75, 2 => 9276, 3 => 29656, 4 => 4543, 5 => 30699, 6 => 20646, 7 => 21921, 8 => 28050),
    22 => integer_vector_t'(0 => 8, 1 => 76, 2 => 15975, 3 => 25634, 4 => 5520, 5 => 31119, 6 => 13715, 7 => 21949, 8 => 19605),
    23 => integer_vector_t'(0 => 8, 1 => 77, 2 => 18688, 3 => 4608, 4 => 31755, 5 => 30165, 6 => 13103, 7 => 10706, 8 => 29224),
    24 => integer_vector_t'(0 => 8, 1 => 78, 2 => 21514, 3 => 23117, 4 => 12245, 5 => 26035, 6 => 31656, 7 => 25631, 8 => 30699),
    25 => integer_vector_t'(0 => 8, 1 => 79, 2 => 9674, 3 => 24966, 4 => 31285, 5 => 29908, 6 => 17042, 7 => 24588, 8 => 31857),
    26 => integer_vector_t'(0 => 8, 1 => 80, 2 => 21856, 3 => 27777, 4 => 29919, 5 => 27000, 6 => 14897, 7 => 11409, 8 => 7122),
    27 => integer_vector_t'(0 => 8, 1 => 81, 2 => 29773, 3 => 23310, 4 => 263, 5 => 4877, 6 => 28622, 7 => 20545, 8 => 22092),
    28 => integer_vector_t'(0 => 8, 1 => 82, 2 => 15605, 3 => 5651, 4 => 21864, 5 => 3967, 6 => 14419, 7 => 22757, 8 => 15896),
    29 => integer_vector_t'(0 => 8, 1 => 83, 2 => 30145, 3 => 1759, 4 => 10139, 5 => 29223, 6 => 26086, 7 => 10556, 8 => 5098),
    30 => integer_vector_t'(0 => 8, 1 => 84, 2 => 18815, 3 => 16575, 4 => 2936, 5 => 24457, 6 => 26738, 7 => 6030, 8 => 505),
    31 => integer_vector_t'(0 => 8, 1 => 85, 2 => 30326, 3 => 22298, 4 => 27562, 5 => 20131, 6 => 26390, 7 => 6247, 8 => 24791),
    32 => integer_vector_t'(0 => 8, 1 => 86, 2 => 928, 3 => 29246, 4 => 21246, 5 => 12400, 6 => 15311, 7 => 32309, 8 => 18608),
    33 => integer_vector_t'(0 => 8, 1 => 87, 2 => 20314, 3 => 6025, 4 => 26689, 5 => 16302, 6 => 2296, 7 => 3244, 8 => 19613),
    34 => integer_vector_t'(0 => 8, 1 => 88, 2 => 6237, 3 => 11943, 4 => 22851, 5 => 15642, 6 => 23857, 7 => 15112, 8 => 20947),
    35 => integer_vector_t'(0 => 8, 1 => 89, 2 => 26403, 3 => 25168, 4 => 19038, 5 => 18384, 6 => 8882, 7 => 12719, 8 => 7093),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 14567, 3 => 24965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3908, 3 => 100, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10279, 3 => 240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 24102, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 12383, 3 => 4173, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 13861, 3 => 15918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 21327, 3 => 1046, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5288, 3 => 14579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 28158, 3 => 8069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 16583, 3 => 11098, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 16681, 3 => 28363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 13980, 3 => 24725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 32169, 3 => 17989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 10907, 3 => 2767, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 21557, 3 => 3818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 26676, 3 => 12422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 7676, 3 => 8754, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 14905, 3 => 20232, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 15719, 3 => 24646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 31942, 3 => 8589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 19978, 3 => 27197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 27060, 3 => 15071, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6071, 3 => 26649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10393, 3 => 11176, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 9597, 3 => 13370, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7081, 3 => 17677, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 1433, 3 => 19513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 26925, 3 => 9014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 19202, 3 => 8900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 18152, 3 => 30647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20803, 3 => 1737, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 11804, 3 => 25221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 31683, 3 => 17783, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 29694, 3 => 9345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 12280, 3 => 26611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 6526, 3 => 26122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 26165, 3 => 11241, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 7666, 3 => 26962, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 16290, 3 => 8480, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 11774, 3 => 10120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 30051, 3 => 30426, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 1335, 3 => 15424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6865, 3 => 17742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 31779, 3 => 12489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 32120, 3 => 21001, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 14508, 3 => 6996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 979, 3 => 25024, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 4554, 3 => 21896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 7989, 3 => 21777, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 4972, 3 => 20661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 6612, 3 => 2730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 12742, 3 => 4418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 29194, 3 => 595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 19267, 3 => 20113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_3.csv, table is 60x196 (1470.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3 : integer_2d_array_t(0 to 59)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 34903, 2 => 20927, 3 => 32093, 4 => 1052, 5 => 25611, 6 => 16093, 7 => 16454, 8 => 5520, 9 => 506, 10 => 37399, 11 => 18518, 12 => 21120),
    1 => integer_vector_t'(0 => 12, 1 => 11636, 2 => 14594, 3 => 22158, 4 => 14763, 5 => 15333, 6 => 6838, 7 => 22222, 8 => 37856, 9 => 14985, 10 => 31041, 11 => 18704, 12 => 32910),
    2 => integer_vector_t'(0 => 12, 1 => 17449, 2 => 1665, 3 => 35639, 4 => 16624, 5 => 12867, 6 => 12449, 7 => 10241, 8 => 11650, 9 => 25622, 10 => 34372, 11 => 19878, 12 => 26894),
    3 => integer_vector_t'(0 => 12, 1 => 29235, 2 => 19780, 3 => 36056, 4 => 20129, 5 => 20029, 6 => 5457, 7 => 8157, 8 => 35554, 9 => 21237, 10 => 7943, 11 => 13873, 12 => 14980),
    4 => integer_vector_t'(0 => 12, 1 => 9912, 2 => 7143, 3 => 35911, 4 => 12043, 5 => 17360, 6 => 37253, 7 => 25588, 8 => 11827, 9 => 29152, 10 => 21936, 11 => 24125, 12 => 40870),
    5 => integer_vector_t'(0 => 12, 1 => 40701, 2 => 36035, 3 => 39556, 4 => 12366, 5 => 19946, 6 => 29072, 7 => 16365, 8 => 35495, 9 => 22686, 10 => 11106, 11 => 8756, 12 => 34863),
    6 => integer_vector_t'(0 => 12, 1 => 19165, 2 => 15702, 3 => 13536, 4 => 40238, 5 => 4465, 6 => 40034, 7 => 40590, 8 => 37540, 9 => 17162, 10 => 1712, 11 => 20577, 12 => 14138),
    7 => integer_vector_t'(0 => 12, 1 => 31338, 2 => 19342, 3 => 9301, 4 => 39375, 5 => 3211, 6 => 1316, 7 => 33409, 8 => 28670, 9 => 12282, 10 => 6118, 11 => 29236, 12 => 35787),
    8 => integer_vector_t'(0 => 12, 1 => 11504, 2 => 30506, 3 => 19558, 4 => 5100, 5 => 24188, 6 => 24738, 7 => 30397, 8 => 33775, 9 => 9699, 10 => 6215, 11 => 3397, 12 => 37451),
    9 => integer_vector_t'(0 => 12, 1 => 34689, 2 => 23126, 3 => 7571, 4 => 1058, 5 => 12127, 6 => 27518, 7 => 23064, 8 => 11265, 9 => 14867, 10 => 30451, 11 => 28289, 12 => 2966),
    10 => integer_vector_t'(0 => 12, 1 => 11660, 2 => 15334, 3 => 16867, 4 => 15160, 5 => 38343, 6 => 3778, 7 => 4265, 8 => 39139, 9 => 17293, 10 => 26229, 11 => 42604, 12 => 13486),
    11 => integer_vector_t'(0 => 12, 1 => 31497, 2 => 1365, 3 => 14828, 4 => 7453, 5 => 26350, 6 => 41346, 7 => 28643, 8 => 23421, 9 => 8354, 10 => 16255, 11 => 11055, 12 => 24279),
    12 => integer_vector_t'(0 => 12, 1 => 15687, 2 => 12467, 3 => 13906, 4 => 5215, 5 => 41328, 6 => 23755, 7 => 20800, 8 => 6447, 9 => 7970, 10 => 2803, 11 => 33262, 12 => 39843),
    13 => integer_vector_t'(0 => 12, 1 => 5363, 2 => 22469, 3 => 38091, 4 => 28457, 5 => 36696, 6 => 34471, 7 => 23619, 8 => 2404, 9 => 24229, 10 => 41754, 11 => 1297, 12 => 18563),
    14 => integer_vector_t'(0 => 12, 1 => 3673, 2 => 39070, 3 => 14480, 4 => 30279, 5 => 37483, 6 => 7580, 7 => 29519, 8 => 30519, 9 => 39831, 10 => 20252, 11 => 18132, 12 => 20010),
    15 => integer_vector_t'(0 => 12, 1 => 34386, 2 => 7252, 3 => 27526, 4 => 12950, 5 => 6875, 6 => 43020, 7 => 31566, 8 => 39069, 9 => 18985, 10 => 15541, 11 => 40020, 12 => 16715),
    16 => integer_vector_t'(0 => 12, 1 => 1721, 2 => 37332, 3 => 39953, 4 => 17430, 5 => 32134, 6 => 29162, 7 => 10490, 8 => 12971, 9 => 28581, 10 => 29331, 11 => 6489, 12 => 35383),
    17 => integer_vector_t'(0 => 12, 1 => 736, 2 => 7022, 3 => 42349, 4 => 8783, 5 => 6767, 6 => 11871, 7 => 21675, 8 => 10325, 9 => 11548, 10 => 25978, 11 => 431, 12 => 24085),
    18 => integer_vector_t'(0 => 12, 1 => 1925, 2 => 10602, 3 => 28585, 4 => 12170, 5 => 15156, 6 => 34404, 7 => 8351, 8 => 13273, 9 => 20208, 10 => 5800, 11 => 15367, 12 => 21764),
    19 => integer_vector_t'(0 => 12, 1 => 16279, 2 => 37832, 3 => 34792, 4 => 21250, 5 => 34192, 6 => 7406, 7 => 41488, 8 => 18346, 9 => 29227, 10 => 26127, 11 => 25493, 12 => 7048),
    20 => integer_vector_t'(0 => 3, 1 => 39948, 2 => 28229, 3 => 24899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 17408, 2 => 14274, 3 => 38993, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 38774, 2 => 15968, 3 => 28459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 41404, 2 => 27249, 3 => 27425, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 41229, 2 => 6082, 3 => 43114, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 13957, 2 => 4979, 3 => 40654, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 3093, 2 => 3438, 3 => 34992, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 34082, 2 => 6172, 3 => 28760, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 42210, 2 => 34141, 3 => 41021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14705, 2 => 17783, 3 => 10134, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 41755, 2 => 39884, 3 => 22773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14615, 2 => 15593, 3 => 1642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 29111, 2 => 37061, 3 => 39860, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 9579, 2 => 33552, 3 => 633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 12951, 2 => 21137, 3 => 39608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 38244, 2 => 27361, 3 => 29417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 2939, 2 => 10172, 3 => 36479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 29094, 2 => 5357, 3 => 19224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 9562, 2 => 24436, 3 => 28637, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 40177, 2 => 2326, 3 => 13504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 6834, 2 => 21583, 3 => 42516, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 40651, 2 => 42810, 3 => 25709, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 31557, 2 => 32138, 3 => 38142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 18624, 2 => 41867, 3 => 39296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 37560, 2 => 14295, 3 => 16245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 6821, 2 => 21679, 3 => 31570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 25339, 2 => 25083, 3 => 22081, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 8047, 2 => 697, 3 => 35268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 9884, 2 => 17073, 3 => 19995, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 26848, 2 => 35245, 3 => 8390, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 18658, 2 => 16134, 3 => 14807, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 12201, 2 => 32944, 3 => 5035, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 25236, 2 => 1216, 3 => 38986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 42994, 2 => 24782, 3 => 8681, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 28321, 2 => 4932, 3 => 34249, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 4107, 2 => 29382, 3 => 32124, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 22157, 2 => 2624, 3 => 14468, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 38788, 2 => 27081, 3 => 7936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4368, 2 => 26148, 3 => 10578, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 25353, 2 => 4122, 3 => 39751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_4.csv, table is 45x196 (1102.5 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4 : integer_2d_array_t(0 to 44)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 23606, 2 => 36098, 3 => 1140, 4 => 28859, 5 => 18148, 6 => 18510, 7 => 6226, 8 => 540, 9 => 42014, 10 => 20879, 11 => 23802, 12 => 47088),
    1 => integer_vector_t'(0 => 12, 1 => 16419, 2 => 24928, 3 => 16609, 4 => 17248, 5 => 7693, 6 => 24997, 7 => 42587, 8 => 16858, 9 => 34921, 10 => 21042, 11 => 37024, 12 => 20692),
    2 => integer_vector_t'(0 => 12, 1 => 1874, 2 => 40094, 3 => 18704, 4 => 14474, 5 => 14004, 6 => 11519, 7 => 13106, 8 => 28826, 9 => 38669, 10 => 22363, 11 => 30255, 12 => 31105),
    3 => integer_vector_t'(0 => 12, 1 => 22254, 2 => 40564, 3 => 22645, 4 => 22532, 5 => 6134, 6 => 9176, 7 => 39998, 8 => 23892, 9 => 8937, 10 => 15608, 11 => 16854, 12 => 31009),
    4 => integer_vector_t'(0 => 12, 1 => 8037, 2 => 40401, 3 => 13550, 4 => 19526, 5 => 41902, 6 => 28782, 7 => 13304, 8 => 32796, 9 => 24679, 10 => 27140, 11 => 45980, 12 => 10021),
    5 => integer_vector_t'(0 => 12, 1 => 40540, 2 => 44498, 3 => 13911, 4 => 22435, 5 => 32701, 6 => 18405, 7 => 39929, 8 => 25521, 9 => 12497, 10 => 9851, 11 => 39223, 12 => 34823),
    6 => integer_vector_t'(0 => 12, 1 => 15233, 2 => 45333, 3 => 5041, 4 => 44979, 5 => 45710, 6 => 42150, 7 => 19416, 8 => 1892, 9 => 23121, 10 => 15860, 11 => 8832, 12 => 10308),
    7 => integer_vector_t'(0 => 12, 1 => 10468, 2 => 44296, 3 => 3611, 4 => 1480, 5 => 37581, 6 => 32254, 7 => 13817, 8 => 6883, 9 => 32892, 10 => 40258, 11 => 46538, 12 => 11940),
    8 => integer_vector_t'(0 => 12, 1 => 6705, 2 => 21634, 3 => 28150, 4 => 43757, 5 => 895, 6 => 6547, 7 => 20970, 8 => 28914, 9 => 30117, 10 => 25736, 11 => 41734, 12 => 11392),
    9 => integer_vector_t'(0 => 12, 1 => 22002, 2 => 5739, 3 => 27210, 4 => 27828, 5 => 34192, 6 => 37992, 7 => 10915, 8 => 6998, 9 => 3824, 10 => 42130, 11 => 4494, 12 => 35739),
    10 => integer_vector_t'(0 => 12, 1 => 8515, 2 => 1191, 3 => 13642, 4 => 30950, 5 => 25943, 6 => 12673, 7 => 16726, 8 => 34261, 9 => 31828, 10 => 3340, 11 => 8747, 12 => 39225),
    11 => integer_vector_t'(0 => 12, 1 => 18979, 2 => 17058, 3 => 43130, 4 => 4246, 5 => 4793, 6 => 44030, 7 => 19454, 8 => 29511, 9 => 47929, 10 => 15174, 11 => 24333, 12 => 19354),
    12 => integer_vector_t'(0 => 12, 1 => 16694, 2 => 8381, 3 => 29642, 4 => 46516, 5 => 32224, 6 => 26344, 7 => 9405, 8 => 18292, 9 => 12437, 10 => 27316, 11 => 35466, 12 => 41992),
    13 => integer_vector_t'(0 => 12, 1 => 15642, 2 => 5871, 3 => 46489, 4 => 26723, 5 => 23396, 6 => 7257, 7 => 8974, 8 => 3156, 9 => 37420, 10 => 44823, 11 => 35423, 12 => 13541),
    14 => integer_vector_t'(0 => 12, 1 => 42858, 2 => 32008, 3 => 41282, 4 => 38773, 5 => 26570, 6 => 2702, 7 => 27260, 8 => 46974, 9 => 1469, 10 => 20887, 11 => 27426, 12 => 38553),
    15 => integer_vector_t'(0 => 3, 1 => 22152, 2 => 24261, 3 => 8297, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 19347, 2 => 9978, 3 => 27802, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 34991, 2 => 6354, 3 => 33561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 29782, 2 => 30875, 3 => 29523, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 9278, 2 => 48512, 3 => 14349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 38061, 2 => 4165, 3 => 43878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 8548, 2 => 33172, 3 => 34410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22535, 2 => 28811, 3 => 23950, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 20439, 2 => 4027, 3 => 24186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 38618, 2 => 8187, 3 => 30947, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 35538, 2 => 43880, 3 => 21459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 7091, 2 => 45616, 3 => 15063, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 5505, 2 => 9315, 3 => 21908, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 36046, 2 => 32914, 3 => 11836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 7304, 2 => 39782, 3 => 33721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 16905, 2 => 29962, 3 => 12980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11171, 2 => 23709, 3 => 22460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 34541, 2 => 9937, 3 => 44500, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 14035, 2 => 47316, 3 => 8815, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 15057, 2 => 45482, 3 => 24461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 30518, 2 => 36877, 3 => 879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7583, 2 => 13364, 3 => 24332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 448, 2 => 27056, 3 => 4682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 12083, 2 => 31378, 3 => 21670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 1159, 2 => 18031, 3 => 2221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 17028, 2 => 38715, 3 => 9350, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 17343, 2 => 24530, 3 => 29574, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 46128, 2 => 31039, 3 => 32818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 20373, 2 => 36967, 3 => 18345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 46685, 2 => 20622, 3 => 32806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_3.csv, table is 120x189 (2835.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 14, 9 => 15, 10 => 15, 11 => 15, 12 => 15, 13 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3 : integer_2d_array_t(0 to 119)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 10491, 3 => 16043, 4 => 506, 5 => 12826, 6 => 8065, 7 => 8226, 8 => 2767, 9 => 240, 10 => 18673, 11 => 9279, 12 => 10579, 13 => 20928),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 17819, 3 => 8313, 4 => 6433, 5 => 6224, 6 => 5120, 7 => 5824, 8 => 12812, 9 => 17187, 10 => 9940, 11 => 13447, 12 => 13825, 13 => 18483),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 17957, 3 => 6024, 4 => 8681, 5 => 18628, 6 => 12794, 7 => 5915, 8 => 14576, 9 => 10970, 10 => 12064, 11 => 20437, 12 => 4455, 13 => 7151),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 19777, 3 => 6183, 4 => 9972, 5 => 14536, 6 => 8182, 7 => 17749, 8 => 11341, 9 => 5556, 10 => 4379, 11 => 17434, 12 => 15477, 13 => 18532),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 4651, 3 => 19689, 4 => 1608, 5 => 659, 6 => 16707, 7 => 14335, 8 => 6143, 9 => 3058, 10 => 14618, 11 => 17894, 12 => 20684, 13 => 5306),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 9778, 3 => 2552, 4 => 12096, 5 => 12369, 6 => 15198, 7 => 16890, 8 => 4851, 9 => 3109, 10 => 1700, 11 => 18725, 12 => 1997, 13 => 15882),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 486, 3 => 6111, 4 => 13743, 5 => 11537, 6 => 5591, 7 => 7433, 8 => 15227, 9 => 14145, 10 => 1483, 11 => 3887, 12 => 17431, 13 => 12430),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 20647, 3 => 14311, 4 => 11734, 5 => 4180, 6 => 8110, 7 => 5525, 8 => 12141, 9 => 15761, 10 => 18661, 11 => 18441, 12 => 10569, 13 => 8192),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 3791, 3 => 14759, 4 => 15264, 5 => 19918, 6 => 10132, 7 => 9062, 8 => 10010, 9 => 12786, 10 => 10675, 11 => 9682, 12 => 19246, 13 => 5454),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 19525, 3 => 9485, 4 => 7777, 5 => 19999, 6 => 8378, 7 => 9209, 8 => 3163, 9 => 20232, 10 => 6690, 11 => 16518, 12 => 716, 13 => 7353),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 4588, 3 => 6709, 4 => 20202, 5 => 10905, 6 => 915, 7 => 4317, 8 => 11073, 9 => 13576, 10 => 16433, 11 => 368, 12 => 3508, 13 => 21171),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 14072, 3 => 4033, 4 => 19959, 5 => 12608, 6 => 631, 7 => 19494, 8 => 14160, 9 => 8249, 10 => 10223, 11 => 21504, 12 => 12395, 13 => 4322),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 13800, 3 => 14161, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2948, 3 => 9647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 14693, 3 => 16027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 20506, 3 => 11082, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1143, 3 => 9020, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13501, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1548, 3 => 2190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 12216, 3 => 21556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 19897, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4189, 3 => 7958, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 15940, 3 => 10048, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 515, 3 => 12614, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8501, 3 => 8450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 17595, 3 => 16784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 5913, 3 => 8495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 16394, 3 => 10423, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7409, 3 => 6981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6678, 3 => 15939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20344, 3 => 12987, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 2510, 3 => 14588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 17918, 3 => 6655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 6703, 3 => 19451, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 496, 3 => 4217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7290, 3 => 5766, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 10521, 3 => 8925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 20379, 3 => 11905, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4090, 3 => 5838, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 19082, 3 => 17040, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 20233, 3 => 12352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 19365, 3 => 19546, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6249, 3 => 19030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11037, 3 => 19193, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 19760, 3 => 11772, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 45, 2 => 19644, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16076, 3 => 3521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11779, 3 => 21062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 48, 2 => 13062, 3 => 9682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 49, 2 => 8934, 3 => 5217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 50, 2 => 11087, 3 => 3319, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 51, 2 => 18892, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 52, 2 => 7894, 3 => 3898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 53, 2 => 5963, 3 => 4360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 54, 2 => 7346, 3 => 11726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5182, 3 => 5609, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 56, 2 => 2412, 3 => 17295, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 57, 2 => 9845, 3 => 20494, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 58, 2 => 6687, 3 => 1864, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 59, 2 => 20564, 3 => 5216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18226, 3 => 17207, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9380, 3 => 8266, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7073, 3 => 3065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 18252, 3 => 13437, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9161, 3 => 15642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10714, 3 => 10153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 11585, 3 => 9078, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5359, 3 => 9418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 9024, 3 => 9515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1206, 3 => 16354, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 14994, 3 => 1102, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9375, 3 => 20796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 15964, 3 => 6027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14789, 3 => 6452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8002, 3 => 18591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 14742, 3 => 14089, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 253, 3 => 3045, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1274, 3 => 19286, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 14777, 3 => 2044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 13920, 3 => 9900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 452, 3 => 7374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 18206, 3 => 9921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6131, 3 => 5414, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10077, 3 => 9726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 12045, 3 => 5479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4322, 3 => 7990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 15616, 3 => 5550, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 15561, 3 => 10661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 20718, 3 => 7387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2518, 3 => 18804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8984, 3 => 2600, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6516, 3 => 17909, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 32, 2 => 11148, 3 => 98, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 33, 2 => 20559, 3 => 3704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7510, 3 => 1569, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 35, 2 => 16000, 3 => 11692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 36, 2 => 9147, 3 => 10303, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 37, 2 => 16650, 3 => 191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15577, 3 => 18685, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 39, 2 => 17167, 3 => 20917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 40, 2 => 4256, 3 => 3391, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 41, 2 => 20092, 3 => 17219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 42, 2 => 9218, 3 => 5056, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 43, 2 => 18429, 3 => 8472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12093, 3 => 20753, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 45, 2 => 16345, 3 => 12748, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16023, 3 => 11095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 47, 2 => 5048, 3 => 17595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 48, 2 => 18995, 3 => 4817, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 49, 2 => 16483, 3 => 3536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 50, 2 => 1439, 3 => 16148, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 51, 2 => 3661, 3 => 3039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 52, 2 => 19010, 3 => 18121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 53, 2 => 8968, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 54, 2 => 13427, 3 => 18003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5303, 3 => 3083, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 56, 2 => 531, 3 => 16668, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 57, 2 => 4771, 3 => 6722, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 58, 2 => 5695, 3 => 7960, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 59, 2 => 3589, 3 => 14630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_5.csv, table is 72x196 (1764.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5 : integer_2d_array_t(0 to 71)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 31413, 2 => 18834, 3 => 28884, 4 => 947, 5 => 23050, 6 => 14484, 7 => 14809, 8 => 4968, 9 => 455, 10 => 33659, 11 => 16666, 12 => 19008),
    1 => integer_vector_t'(0 => 12, 1 => 13172, 2 => 19939, 3 => 13354, 4 => 13719, 5 => 6132, 6 => 20086, 7 => 34040, 8 => 13442, 9 => 27958, 10 => 16813, 11 => 29619, 12 => 16553),
    2 => integer_vector_t'(0 => 12, 1 => 1499, 2 => 32075, 3 => 14962, 4 => 11578, 5 => 11204, 6 => 9217, 7 => 10485, 8 => 23062, 9 => 30936, 10 => 17892, 11 => 24204, 12 => 24885),
    3 => integer_vector_t'(0 => 12, 1 => 32490, 2 => 18086, 3 => 18007, 4 => 4957, 5 => 7285, 6 => 32073, 7 => 19038, 8 => 7152, 9 => 12486, 10 => 13483, 11 => 24808, 12 => 21759),
    4 => integer_vector_t'(0 => 12, 1 => 32321, 2 => 10839, 3 => 15620, 4 => 33521, 5 => 23030, 6 => 10646, 7 => 26236, 8 => 19744, 9 => 21713, 10 => 36784, 11 => 8016, 12 => 12869),
    5 => integer_vector_t'(0 => 12, 1 => 35597, 2 => 11129, 3 => 17948, 4 => 26160, 5 => 14729, 6 => 31943, 7 => 20416, 8 => 10000, 9 => 7882, 10 => 31380, 11 => 27858, 12 => 33356),
    6 => integer_vector_t'(0 => 12, 1 => 14125, 2 => 12131, 3 => 36199, 4 => 4058, 5 => 35992, 6 => 36594, 7 => 33698, 8 => 15475, 9 => 1566, 10 => 18498, 11 => 12725, 12 => 7067),
    7 => integer_vector_t'(0 => 12, 1 => 17406, 2 => 8372, 3 => 35437, 4 => 2888, 5 => 1184, 6 => 30068, 7 => 25802, 8 => 11056, 9 => 5507, 10 => 26313, 11 => 32205, 12 => 37232),
    8 => integer_vector_t'(0 => 12, 1 => 15254, 2 => 5365, 3 => 17308, 4 => 22519, 5 => 35009, 6 => 718, 7 => 5240, 8 => 16778, 9 => 23131, 10 => 24092, 11 => 20587, 12 => 33385),
    9 => integer_vector_t'(0 => 12, 1 => 27455, 2 => 17602, 3 => 4590, 4 => 21767, 5 => 22266, 6 => 27357, 7 => 30400, 8 => 8732, 9 => 5596, 10 => 3060, 11 => 33703, 12 => 3596),
    10 => integer_vector_t'(0 => 12, 1 => 6882, 2 => 873, 3 => 10997, 4 => 24738, 5 => 20770, 6 => 10067, 7 => 13379, 8 => 27409, 9 => 25463, 10 => 2673, 11 => 6998, 12 => 31378),
    11 => integer_vector_t'(0 => 12, 1 => 15181, 2 => 13645, 3 => 34501, 4 => 3393, 5 => 3840, 6 => 35227, 7 => 15562, 8 => 23615, 9 => 38342, 10 => 12139, 11 => 19471, 12 => 15483),
    12 => integer_vector_t'(0 => 12, 1 => 13350, 2 => 6707, 3 => 23709, 4 => 37204, 5 => 25778, 6 => 21082, 7 => 7511, 8 => 14588, 9 => 10010, 10 => 21854, 11 => 28375, 12 => 33591),
    13 => integer_vector_t'(0 => 12, 1 => 12514, 2 => 4695, 3 => 37190, 4 => 21379, 5 => 18723, 6 => 5802, 7 => 7182, 8 => 2529, 9 => 29936, 10 => 35860, 11 => 28338, 12 => 10835),
    14 => integer_vector_t'(0 => 12, 1 => 34283, 2 => 25610, 3 => 33026, 4 => 31017, 5 => 21259, 6 => 2165, 7 => 21807, 8 => 37578, 9 => 1175, 10 => 16710, 11 => 21939, 12 => 30841),
    15 => integer_vector_t'(0 => 12, 1 => 27292, 2 => 33730, 3 => 6836, 4 => 26476, 5 => 27539, 6 => 35784, 7 => 18245, 8 => 16394, 9 => 17939, 10 => 23094, 11 => 19216, 12 => 17432),
    16 => integer_vector_t'(0 => 12, 1 => 11655, 2 => 6183, 3 => 38708, 4 => 28408, 5 => 35157, 6 => 17089, 7 => 13998, 8 => 36029, 9 => 15052, 10 => 16617, 11 => 5638, 12 => 36464),
    17 => integer_vector_t'(0 => 12, 1 => 15693, 2 => 28923, 3 => 26245, 4 => 9432, 5 => 11675, 6 => 25720, 7 => 26405, 8 => 5838, 9 => 31851, 10 => 26898, 11 => 8090, 12 => 37037),
    18 => integer_vector_t'(0 => 12, 1 => 24418, 2 => 27583, 3 => 7959, 4 => 35562, 5 => 37771, 6 => 17784, 7 => 11382, 8 => 11156, 9 => 37855, 10 => 7073, 11 => 21685, 12 => 34515),
    19 => integer_vector_t'(0 => 12, 1 => 10977, 2 => 13633, 3 => 30969, 4 => 7516, 5 => 11943, 6 => 18199, 7 => 5231, 8 => 13825, 9 => 19589, 10 => 23661, 11 => 11150, 12 => 35602),
    20 => integer_vector_t'(0 => 12, 1 => 19124, 2 => 30774, 3 => 6670, 4 => 37344, 5 => 16510, 6 => 26317, 7 => 23518, 8 => 22957, 9 => 6348, 10 => 34069, 11 => 8845, 12 => 20175),
    21 => integer_vector_t'(0 => 12, 1 => 34985, 2 => 14441, 3 => 25668, 4 => 4116, 5 => 3019, 6 => 21049, 7 => 37308, 8 => 24551, 9 => 24727, 10 => 20104, 11 => 24850, 12 => 12114),
    22 => integer_vector_t'(0 => 12, 1 => 38187, 2 => 28527, 3 => 13108, 4 => 13985, 5 => 1425, 6 => 21477, 7 => 30807, 8 => 8613, 9 => 26241, 10 => 33368, 11 => 35913, 12 => 32477),
    23 => integer_vector_t'(0 => 12, 1 => 5903, 2 => 34390, 3 => 24641, 4 => 26556, 5 => 23007, 6 => 27305, 7 => 38247, 8 => 2621, 9 => 9122, 10 => 32806, 11 => 21554, 12 => 18685),
    24 => integer_vector_t'(0 => 3, 1 => 17287, 2 => 27292, 3 => 19033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25796, 2 => 31795, 3 => 12152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 12184, 2 => 35088, 3 => 31226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 38263, 2 => 33386, 3 => 24892, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 23114, 2 => 37995, 3 => 29796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 34336, 2 => 10551, 3 => 36245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 35407, 2 => 175, 3 => 7203, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14654, 2 => 38201, 3 => 22605, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 28404, 2 => 6595, 3 => 1018, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 19932, 2 => 3524, 3 => 29305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 31749, 2 => 20247, 3 => 8128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 18026, 2 => 36357, 3 => 26735, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7543, 2 => 29767, 3 => 13588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 13333, 2 => 25965, 3 => 8463, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 14504, 2 => 36796, 3 => 19710, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4528, 2 => 25299, 3 => 7318, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 35091, 2 => 25550, 3 => 14798, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 7824, 2 => 215, 3 => 1248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 30848, 2 => 5362, 3 => 17291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 28932, 2 => 30249, 3 => 27073, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 13062, 2 => 2103, 3 => 16206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 7129, 2 => 32062, 3 => 19612, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 9512, 2 => 21936, 3 => 38833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 35849, 2 => 33754, 3 => 23450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18705, 2 => 28656, 3 => 18111, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 22749, 2 => 27456, 3 => 32187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 28229, 2 => 31684, 3 => 30160, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15293, 2 => 8483, 3 => 28002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 14880, 2 => 13334, 3 => 12584, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 28646, 2 => 2558, 3 => 19687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 6259, 2 => 4499, 3 => 26336, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 11952, 2 => 28386, 3 => 8405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 10609, 2 => 961, 3 => 7582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 10423, 2 => 13191, 3 => 26818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 15922, 2 => 36654, 3 => 21450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 10492, 2 => 1532, 3 => 1205, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 30551, 2 => 36482, 3 => 22153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 5156, 2 => 11330, 3 => 34243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 28616, 2 => 35369, 3 => 13322, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 8962, 2 => 1485, 3 => 21186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 23541, 2 => 17445, 3 => 35561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 33133, 2 => 11593, 3 => 19895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 33917, 2 => 7863, 3 => 33651, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 20063, 2 => 28331, 3 => 10702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 13195, 2 => 21107, 3 => 21859, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 4364, 2 => 31137, 3 => 4804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 5585, 2 => 2037, 3 => 4830, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 30672, 2 => 16927, 3 => 14800, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_4.csv, table is 135x164 (2767.5 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4 : integer_2d_array_t(0 to 134)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 0, 2 => 6385, 3 => 7901, 4 => 14611, 5 => 13389, 6 => 11200, 7 => 3252, 8 => 5243, 9 => 2504, 10 => 2722, 11 => 821, 12 => 7374),
    1 => integer_vector_t'(0 => 12, 1 => 1, 2 => 11359, 3 => 2698, 4 => 357, 5 => 13824, 6 => 12772, 7 => 7244, 8 => 6752, 9 => 15310, 10 => 852, 11 => 2001, 12 => 11417),
    2 => integer_vector_t'(0 => 12, 1 => 2, 2 => 7862, 3 => 7977, 4 => 6321, 5 => 13612, 6 => 12197, 7 => 14449, 8 => 15137, 9 => 13860, 10 => 1708, 11 => 6399, 12 => 13444),
    3 => integer_vector_t'(0 => 12, 1 => 3, 2 => 1560, 3 => 11804, 4 => 6975, 5 => 13292, 6 => 3646, 7 => 3812, 8 => 8772, 9 => 7306, 10 => 5795, 11 => 14327, 12 => 7866),
    4 => integer_vector_t'(0 => 12, 1 => 4, 2 => 7626, 3 => 11407, 4 => 14599, 5 => 9689, 6 => 1628, 7 => 2113, 8 => 10809, 9 => 9283, 10 => 1230, 11 => 15241, 12 => 4870),
    5 => integer_vector_t'(0 => 12, 1 => 5, 2 => 1610, 3 => 5699, 4 => 15876, 5 => 9446, 6 => 12515, 7 => 1400, 8 => 6303, 9 => 5411, 10 => 14181, 11 => 13925, 12 => 7358),
    6 => integer_vector_t'(0 => 12, 1 => 6, 2 => 4059, 3 => 8836, 4 => 3405, 5 => 7853, 6 => 7992, 7 => 15336, 8 => 5970, 9 => 10368, 10 => 10278, 11 => 9675, 12 => 4651),
    7 => integer_vector_t'(0 => 12, 1 => 7, 2 => 4441, 3 => 3963, 4 => 9153, 5 => 2109, 6 => 12683, 7 => 7459, 8 => 12030, 9 => 12221, 10 => 629, 11 => 15212, 12 => 406),
    8 => integer_vector_t'(0 => 12, 1 => 8, 2 => 6007, 3 => 8411, 4 => 5771, 5 => 3497, 6 => 543, 7 => 14202, 8 => 875, 9 => 9186, 10 => 6235, 11 => 13908, 12 => 3563),
    9 => integer_vector_t'(0 => 12, 1 => 9, 2 => 3232, 3 => 6625, 4 => 4795, 5 => 546, 6 => 9781, 7 => 2071, 8 => 7312, 9 => 3399, 10 => 7250, 11 => 4932, 12 => 12652),
    10 => integer_vector_t'(0 => 12, 1 => 10, 2 => 8820, 3 => 10088, 4 => 11090, 5 => 7069, 6 => 6585, 7 => 13134, 8 => 10158, 9 => 7183, 10 => 488, 11 => 7455, 12 => 9238),
    11 => integer_vector_t'(0 => 12, 1 => 11, 2 => 1903, 3 => 10818, 4 => 119, 5 => 215, 6 => 7558, 7 => 11046, 8 => 10615, 9 => 11545, 10 => 14784, 11 => 7961, 12 => 15619),
    12 => integer_vector_t'(0 => 12, 1 => 12, 2 => 3655, 3 => 8736, 4 => 4917, 5 => 15874, 6 => 5129, 7 => 2134, 8 => 15944, 9 => 14768, 10 => 7150, 11 => 2692, 12 => 1469),
    13 => integer_vector_t'(0 => 12, 1 => 13, 2 => 8316, 3 => 3820, 4 => 505, 5 => 8923, 6 => 6757, 7 => 806, 8 => 7957, 9 => 4216, 10 => 15589, 11 => 13244, 12 => 2622),
    14 => integer_vector_t'(0 => 12, 1 => 14, 2 => 14463, 3 => 4852, 4 => 15733, 5 => 3041, 6 => 11193, 7 => 12860, 8 => 13673, 9 => 8152, 10 => 6551, 11 => 15108, 12 => 8758),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3149, 3 => 11981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 13416, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13098, 3 => 13352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 2009, 3 => 14460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 7207, 3 => 4314, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 3312, 3 => 3945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4418, 3 => 6248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 2669, 3 => 13975, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 7571, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14172, 3 => 2967, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7271, 3 => 7138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6135, 3 => 13670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 7490, 3 => 14559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8657, 3 => 2466, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8599, 3 => 12834, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 3470, 3 => 3152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13917, 3 => 4365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 6024, 3 => 13730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 10973, 3 => 14182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 2464, 3 => 13167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 5281, 3 => 15049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 1103, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 2058, 3 => 1069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 9654, 3 => 6095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 14311, 3 => 7667, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 15617, 3 => 8146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 4588, 3 => 11218, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 13660, 3 => 6243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 8578, 3 => 7874, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 11741, 3 => 2686, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1022, 3 => 1264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 1, 2 => 12604, 3 => 9965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 2, 2 => 8217, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3156, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 4, 2 => 354, 3 => 1514, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6978, 3 => 14058, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 6, 2 => 7922, 3 => 16079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 7, 2 => 15087, 3 => 12138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5053, 3 => 6470, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 9, 2 => 12687, 3 => 14932, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15458, 3 => 1763, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8121, 3 => 1721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 12, 2 => 12431, 3 => 549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4129, 3 => 7091, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1426, 3 => 8415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9783, 3 => 7604, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6295, 3 => 11329, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1409, 3 => 12061, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 18, 2 => 8065, 3 => 9087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2918, 3 => 8438, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1293, 3 => 14115, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 21, 2 => 3922, 3 => 13851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3851, 3 => 4000, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5865, 3 => 1768, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2655, 3 => 14957, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 25, 2 => 5565, 3 => 6332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4303, 3 => 12631, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11653, 3 => 12236, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 28, 2 => 16025, 3 => 7632, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4655, 3 => 14128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 30, 2 => 9584, 3 => 13123, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13987, 3 => 9597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 32, 2 => 15409, 3 => 12110, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 33, 2 => 8754, 3 => 15490, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7416, 3 => 15325, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2909, 3 => 15549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 36, 2 => 2995, 3 => 8257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 37, 2 => 9406, 3 => 4791, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 38, 2 => 11111, 3 => 4854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 39, 2 => 2812, 3 => 8521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 40, 2 => 8476, 3 => 14717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7820, 3 => 15360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 42, 2 => 1179, 3 => 7939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 43, 2 => 2357, 3 => 8678, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 44, 2 => 7703, 3 => 6216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3477, 3 => 7067, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3931, 3 => 13845, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7675, 3 => 12899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1754, 3 => 8187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7785, 3 => 1400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 9213, 3 => 5891, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2494, 3 => 7703, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2576, 3 => 7902, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4821, 3 => 15682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 10426, 3 => 11935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1810, 3 => 904, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 11332, 3 => 9264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11312, 3 => 3570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14916, 3 => 2650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7679, 3 => 7842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6089, 3 => 13084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3938, 3 => 2751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8509, 3 => 4648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 12204, 3 => 8917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5749, 3 => 12443, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12613, 3 => 4431, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1344, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 8488, 3 => 13850, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1730, 3 => 14896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14942, 3 => 7126, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 14983, 3 => 8863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6578, 3 => 8564, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 4947, 3 => 396, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 297, 3 => 12805, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 13878, 3 => 6692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11857, 3 => 11186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 31, 2 => 14395, 3 => 11493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 32, 2 => 16145, 3 => 12251, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 33, 2 => 13462, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 34, 2 => 14526, 3 => 13119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2535, 3 => 11243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 36, 2 => 6465, 3 => 12690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 37, 2 => 6872, 3 => 9334, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15371, 3 => 14023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 39, 2 => 8101, 3 => 10187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 40, 2 => 11963, 3 => 4848, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 41, 2 => 15125, 3 => 6119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 42, 2 => 8051, 3 => 14465, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11139, 3 => 5167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 44, 2 => 2883, 3 => 14521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_5.csv, table is 108x184 (2484.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 15, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15, 9 => 15, 10 => 15, 11 => 15, 12 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5 : integer_2d_array_t(0 to 107)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 22422, 2 => 10282, 3 => 11626, 4 => 19997, 5 => 11161, 6 => 2922, 7 => 3122, 8 => 99, 9 => 5625, 10 => 17064, 11 => 8270, 12 => 179),
    1 => integer_vector_t'(0 => 12, 1 => 25087, 2 => 16218, 3 => 17015, 4 => 828, 5 => 20041, 6 => 25656, 7 => 4186, 8 => 11629, 9 => 22599, 10 => 17305, 11 => 22515, 12 => 6463),
    2 => integer_vector_t'(0 => 12, 1 => 11049, 2 => 22853, 3 => 25706, 4 => 14388, 5 => 5500, 6 => 19245, 7 => 8732, 8 => 2177, 9 => 13555, 10 => 11346, 11 => 17265, 12 => 3069),
    3 => integer_vector_t'(0 => 12, 1 => 16581, 2 => 22225, 3 => 12563, 4 => 19717, 5 => 23577, 6 => 11555, 7 => 25496, 8 => 6853, 9 => 25403, 10 => 5218, 11 => 15925, 12 => 21766),
    4 => integer_vector_t'(0 => 12, 1 => 16529, 2 => 14487, 3 => 7643, 4 => 10715, 5 => 17442, 6 => 11119, 7 => 5679, 8 => 14155, 9 => 24213, 10 => 21000, 11 => 1116, 12 => 15620),
    5 => integer_vector_t'(0 => 12, 1 => 5340, 2 => 8636, 3 => 16693, 4 => 1434, 5 => 5635, 6 => 6516, 7 => 9482, 8 => 20189, 9 => 1066, 10 => 15013, 11 => 25361, 12 => 14243),
    6 => integer_vector_t'(0 => 12, 1 => 18506, 2 => 22236, 3 => 20912, 4 => 8952, 5 => 5421, 6 => 15691, 7 => 6126, 8 => 21595, 9 => 500, 10 => 6904, 11 => 13059, 12 => 6802),
    7 => integer_vector_t'(0 => 12, 1 => 8433, 2 => 4694, 3 => 5524, 4 => 14216, 5 => 3685, 6 => 19721, 7 => 25420, 8 => 9937, 9 => 23813, 10 => 9047, 11 => 25651, 12 => 16826),
    8 => integer_vector_t'(0 => 12, 1 => 21500, 2 => 24814, 3 => 6344, 4 => 17382, 5 => 7064, 6 => 13929, 7 => 4004, 8 => 16552, 9 => 12818, 10 => 8720, 11 => 5286, 12 => 2206),
    9 => integer_vector_t'(0 => 12, 1 => 22517, 2 => 2429, 3 => 19065, 4 => 2921, 5 => 21611, 6 => 1873, 7 => 7507, 8 => 5661, 9 => 23006, 10 => 23128, 11 => 20543, 12 => 19777),
    10 => integer_vector_t'(0 => 12, 1 => 1770, 2 => 4636, 3 => 20900, 4 => 14931, 5 => 9247, 6 => 12340, 7 => 11008, 8 => 12966, 9 => 4471, 10 => 2731, 11 => 16445, 12 => 791),
    11 => integer_vector_t'(0 => 12, 1 => 6635, 2 => 14556, 3 => 18865, 4 => 22421, 5 => 22124, 6 => 12697, 7 => 9803, 8 => 25485, 9 => 7744, 10 => 18254, 11 => 11313, 12 => 9004),
    12 => integer_vector_t'(0 => 12, 1 => 19982, 2 => 23963, 3 => 18912, 4 => 7206, 5 => 12500, 6 => 4382, 7 => 20067, 8 => 6177, 9 => 21007, 10 => 1195, 11 => 23547, 12 => 24837),
    13 => integer_vector_t'(0 => 12, 1 => 756, 2 => 11158, 3 => 14646, 4 => 20534, 5 => 3647, 6 => 17728, 7 => 11676, 8 => 11843, 9 => 12937, 10 => 4402, 11 => 8261, 12 => 22944),
    14 => integer_vector_t'(0 => 12, 1 => 9306, 2 => 24009, 3 => 10012, 4 => 11081, 5 => 3746, 6 => 24325, 7 => 8060, 8 => 19826, 9 => 842, 10 => 8836, 11 => 2898, 12 => 5019),
    15 => integer_vector_t'(0 => 12, 1 => 7575, 2 => 7455, 3 => 25244, 4 => 4736, 5 => 14400, 6 => 22981, 7 => 5543, 8 => 8006, 9 => 24203, 10 => 13053, 11 => 1120, 12 => 5128),
    16 => integer_vector_t'(0 => 12, 1 => 3482, 2 => 9270, 3 => 13059, 4 => 15825, 5 => 7453, 6 => 23747, 7 => 3656, 8 => 24585, 9 => 16542, 10 => 17507, 11 => 22462, 12 => 14670),
    17 => integer_vector_t'(0 => 12, 1 => 15627, 2 => 15290, 3 => 4198, 4 => 22748, 5 => 5842, 6 => 13395, 7 => 23918, 8 => 16985, 9 => 14929, 10 => 3726, 11 => 25350, 12 => 24157),
    18 => integer_vector_t'(0 => 12, 1 => 24896, 2 => 16365, 3 => 16423, 4 => 13461, 5 => 16615, 6 => 8107, 7 => 24741, 8 => 3604, 9 => 25904, 10 => 8716, 11 => 9604, 12 => 20365),
    19 => integer_vector_t'(0 => 12, 1 => 3729, 2 => 17245, 3 => 18448, 4 => 9862, 5 => 20831, 6 => 25326, 7 => 20517, 8 => 24618, 9 => 13282, 10 => 5099, 11 => 14183, 12 => 8804),
    20 => integer_vector_t'(0 => 12, 1 => 16455, 2 => 17646, 3 => 15376, 4 => 18194, 5 => 25528, 6 => 1777, 7 => 6066, 8 => 21855, 9 => 14372, 10 => 12517, 11 => 4488, 12 => 17490),
    21 => integer_vector_t'(0 => 12, 1 => 1400, 2 => 8135, 3 => 23375, 4 => 20879, 5 => 8476, 6 => 4084, 7 => 12936, 8 => 25536, 9 => 22309, 10 => 16582, 11 => 6402, 12 => 24360),
    22 => integer_vector_t'(0 => 12, 1 => 25119, 2 => 23586, 3 => 128, 4 => 4761, 5 => 10443, 6 => 22536, 7 => 8607, 8 => 9752, 9 => 25446, 10 => 15053, 11 => 1856, 12 => 4040),
    23 => integer_vector_t'(0 => 12, 1 => 377, 2 => 21160, 3 => 13474, 4 => 5451, 5 => 17170, 6 => 5938, 7 => 10256, 8 => 11972, 9 => 24210, 10 => 17833, 11 => 22047, 12 => 16108),
    24 => integer_vector_t'(0 => 12, 1 => 13075, 2 => 9648, 3 => 24546, 4 => 13150, 5 => 23867, 6 => 7309, 7 => 19798, 8 => 2988, 9 => 16858, 10 => 4825, 11 => 23950, 12 => 15125),
    25 => integer_vector_t'(0 => 12, 1 => 20526, 2 => 3553, 3 => 11525, 4 => 23366, 5 => 2452, 6 => 17626, 7 => 19265, 8 => 20172, 9 => 18060, 10 => 24593, 11 => 13255, 12 => 1552),
    26 => integer_vector_t'(0 => 12, 1 => 18839, 2 => 21132, 3 => 20119, 4 => 15214, 5 => 14705, 6 => 7096, 7 => 10174, 8 => 5663, 9 => 18651, 10 => 19700, 11 => 12524, 12 => 14033),
    27 => integer_vector_t'(0 => 12, 1 => 4127, 2 => 2971, 3 => 17499, 4 => 16287, 5 => 22368, 6 => 21463, 7 => 7943, 8 => 18880, 9 => 5567, 10 => 8047, 11 => 23363, 12 => 6797),
    28 => integer_vector_t'(0 => 12, 1 => 10651, 2 => 24471, 3 => 14325, 4 => 4081, 5 => 7258, 6 => 4949, 7 => 7044, 8 => 1078, 9 => 797, 10 => 22910, 11 => 20474, 12 => 4318),
    29 => integer_vector_t'(0 => 12, 1 => 21374, 2 => 13231, 3 => 22985, 4 => 5056, 5 => 3821, 6 => 23718, 7 => 14178, 8 => 9978, 9 => 19030, 10 => 23594, 11 => 8895, 12 => 25358),
    30 => integer_vector_t'(0 => 12, 1 => 6199, 2 => 22056, 3 => 7749, 4 => 13310, 5 => 3999, 6 => 23697, 7 => 16445, 8 => 22636, 9 => 5225, 10 => 22437, 11 => 24153, 12 => 9442),
    31 => integer_vector_t'(0 => 12, 1 => 7978, 2 => 12177, 3 => 2893, 4 => 20778, 5 => 3175, 6 => 8645, 7 => 11863, 8 => 24623, 9 => 10311, 10 => 25767, 11 => 17057, 12 => 3691),
    32 => integer_vector_t'(0 => 12, 1 => 20473, 2 => 11294, 3 => 9914, 4 => 22815, 5 => 2574, 6 => 8439, 7 => 3699, 8 => 5431, 9 => 24840, 10 => 21908, 11 => 16088, 12 => 18244),
    33 => integer_vector_t'(0 => 12, 1 => 8208, 2 => 5755, 3 => 19059, 4 => 8541, 5 => 24924, 6 => 6454, 7 => 11234, 8 => 10492, 9 => 16406, 10 => 10831, 11 => 11436, 12 => 9649),
    34 => integer_vector_t'(0 => 12, 1 => 16264, 2 => 11275, 3 => 24953, 4 => 2347, 5 => 12667, 6 => 19190, 7 => 7257, 8 => 7174, 9 => 24819, 10 => 2938, 11 => 2522, 12 => 11749),
    35 => integer_vector_t'(0 => 12, 1 => 3627, 2 => 5969, 3 => 13862, 4 => 1538, 5 => 23176, 6 => 6353, 7 => 2855, 8 => 17720, 9 => 2472, 10 => 7428, 11 => 573, 12 => 15036),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18539, 3 => 18661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 10502, 3 => 3002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 9368, 3 => 10761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 12299, 3 => 7828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 15048, 3 => 13362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 18444, 3 => 24640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 20775, 3 => 19175, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 18970, 3 => 10971, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5329, 3 => 19982, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 11296, 3 => 18655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15046, 3 => 20659, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 7300, 3 => 22140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 22029, 3 => 14477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 11129, 3 => 742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 13254, 3 => 13813, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 19234, 3 => 13273, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6079, 3 => 21122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 22782, 3 => 5828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 19775, 3 => 4247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1660, 3 => 19413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4403, 3 => 3649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 13371, 3 => 25851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 22770, 3 => 21784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10757, 3 => 14131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 16071, 3 => 21617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 6393, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 597, 3 => 19968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5743, 3 => 8084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 6770, 3 => 9548, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4285, 3 => 17542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 13568, 3 => 22599, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 1786, 3 => 4617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 23238, 3 => 11648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 19627, 3 => 2030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 13601, 3 => 13458, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 13740, 3 => 17328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 25012, 3 => 13944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 22513, 3 => 6687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4934, 3 => 12587, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 21197, 3 => 5133, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 22705, 3 => 6938, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7534, 3 => 24633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 24400, 3 => 12797, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 21911, 3 => 25712, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12039, 3 => 1140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 24306, 3 => 1021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 14012, 3 => 20747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11265, 3 => 15219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 4670, 3 => 15531, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 9417, 3 => 14359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 2415, 3 => 6504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 24964, 3 => 24690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 14443, 3 => 8816, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 6926, 3 => 1291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 54, 2 => 6209, 3 => 20806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 55, 2 => 13915, 3 => 4079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 56, 2 => 24410, 3 => 13196, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 57, 2 => 13505, 3 => 6117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 58, 2 => 9869, 3 => 8220, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 59, 2 => 1570, 3 => 6044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 60, 2 => 25780, 3 => 17387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 61, 2 => 20671, 3 => 24913, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 62, 2 => 24558, 3 => 20591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 63, 2 => 12402, 3 => 3702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 64, 2 => 8314, 3 => 1357, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 65, 2 => 20071, 3 => 14616, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 66, 2 => 17014, 3 => 3688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 67, 2 => 19837, 3 => 946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 68, 2 => 15195, 3 => 12136, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 69, 2 => 7758, 3 => 22808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 70, 2 => 3564, 3 => 2925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 71, 2 => 3434, 3 => 7769, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C4_5.csv, table is 144x150 (2700.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5 : integer_2d_array_t(0 to 143)(0 to 11) := (
    0 => integer_vector_t'(0 => 11, 1 => 0, 2 => 149, 3 => 11212, 4 => 5575, 5 => 6360, 6 => 12559, 7 => 8108, 8 => 8505, 9 => 408, 10 => 10026, 11 => 12828),
    1 => integer_vector_t'(0 => 11, 1 => 1, 2 => 5237, 3 => 490, 4 => 10677, 5 => 4998, 6 => 3869, 7 => 3734, 8 => 3092, 9 => 3509, 10 => 7703, 11 => 10305),
    2 => integer_vector_t'(0 => 11, 1 => 2, 2 => 8742, 3 => 5553, 4 => 2820, 5 => 7085, 6 => 12116, 7 => 10485, 8 => 564, 9 => 7795, 10 => 2972, 11 => 2157),
    3 => integer_vector_t'(0 => 11, 1 => 3, 2 => 2699, 3 => 4304, 4 => 8350, 5 => 712, 6 => 2841, 7 => 3250, 8 => 4731, 9 => 10105, 10 => 517, 11 => 7516),
    4 => integer_vector_t'(0 => 11, 1 => 4, 2 => 12067, 3 => 1351, 4 => 11992, 5 => 12191, 6 => 11267, 7 => 5161, 8 => 537, 9 => 6166, 10 => 4246, 11 => 2363),
    5 => integer_vector_t'(0 => 11, 1 => 5, 2 => 6828, 3 => 7107, 4 => 2127, 5 => 3724, 6 => 5743, 7 => 11040, 8 => 10756, 9 => 4073, 10 => 1011, 11 => 3422),
    6 => integer_vector_t'(0 => 11, 1 => 6, 2 => 11259, 3 => 1216, 4 => 9526, 5 => 1466, 6 => 10816, 7 => 940, 8 => 3744, 9 => 2815, 10 => 11506, 11 => 11573),
    7 => integer_vector_t'(0 => 11, 1 => 7, 2 => 4549, 3 => 11507, 4 => 1118, 5 => 1274, 6 => 11751, 7 => 5207, 8 => 7854, 9 => 12803, 10 => 4047, 11 => 6484),
    8 => integer_vector_t'(0 => 11, 1 => 8, 2 => 8430, 3 => 4115, 4 => 9440, 5 => 413, 6 => 4455, 7 => 2262, 8 => 7915, 9 => 12402, 10 => 8579, 11 => 7052),
    9 => integer_vector_t'(0 => 11, 1 => 9, 2 => 3885, 3 => 9126, 4 => 5665, 5 => 4505, 6 => 2343, 7 => 253, 8 => 4707, 9 => 3742, 10 => 4166, 11 => 1556),
    10 => integer_vector_t'(0 => 11, 1 => 10, 2 => 1704, 3 => 8936, 4 => 6775, 5 => 8639, 6 => 8179, 7 => 7954, 8 => 8234, 9 => 7850, 10 => 8883, 11 => 8713),
    11 => integer_vector_t'(0 => 11, 1 => 11, 2 => 11716, 3 => 4344, 4 => 9087, 5 => 11264, 6 => 2274, 7 => 8832, 8 => 9147, 9 => 11930, 10 => 6054, 11 => 5455),
    12 => integer_vector_t'(0 => 11, 1 => 12, 2 => 7323, 3 => 3970, 4 => 10329, 5 => 2170, 6 => 8262, 7 => 3854, 8 => 2087, 9 => 12899, 10 => 9497, 11 => 11700),
    13 => integer_vector_t'(0 => 11, 1 => 13, 2 => 4418, 3 => 1467, 4 => 2490, 5 => 5841, 6 => 817, 7 => 11453, 8 => 533, 9 => 11217, 10 => 11962, 11 => 5251),
    14 => integer_vector_t'(0 => 11, 1 => 14, 2 => 1541, 3 => 4525, 4 => 7976, 5 => 3457, 6 => 9536, 7 => 7725, 8 => 3788, 9 => 2982, 10 => 6307, 11 => 5997),
    15 => integer_vector_t'(0 => 11, 1 => 15, 2 => 11484, 3 => 2739, 4 => 4023, 5 => 12107, 6 => 6516, 7 => 551, 8 => 2572, 9 => 6628, 10 => 8150, 11 => 9852),
    16 => integer_vector_t'(0 => 11, 1 => 16, 2 => 6070, 3 => 1761, 4 => 4627, 5 => 6534, 6 => 7913, 7 => 3730, 8 => 11866, 9 => 1813, 10 => 12306, 11 => 8249),
    17 => integer_vector_t'(0 => 11, 1 => 17, 2 => 12441, 3 => 5489, 4 => 8748, 5 => 7837, 6 => 7660, 7 => 2102, 8 => 11341, 9 => 2936, 10 => 6712, 11 => 11977),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10155, 3 => 4210, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1010, 3 => 10483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 8900, 3 => 10250, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 10243, 3 => 12278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 7070, 3 => 4397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 12271, 3 => 3887, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 11980, 3 => 6836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 9514, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 7137, 3 => 10281, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11881, 3 => 2526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 1969, 3 => 11477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3044, 3 => 10921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 2236, 3 => 8724, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9104, 3 => 6340, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 7342, 3 => 8582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 11675, 3 => 10405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 6467, 3 => 12775, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 3186, 3 => 12198, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 9621, 3 => 11445, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7486, 3 => 5611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4319, 3 => 4879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2196, 3 => 344, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7527, 3 => 6650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10693, 3 => 2440, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6755, 3 => 2706, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5144, 3 => 5998, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 11043, 3 => 8033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4846, 3 => 4435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4157, 3 => 9228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 12270, 3 => 6562, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11954, 3 => 7592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 7420, 3 => 2592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8810, 3 => 9636, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 689, 3 => 5430, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 920, 3 => 1304, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1253, 3 => 11934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9559, 3 => 6016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 312, 3 => 7589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4439, 3 => 4197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4002, 3 => 9555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12232, 3 => 7779, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1494, 3 => 8782, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 10749, 3 => 3969, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4368, 3 => 3479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6316, 3 => 5342, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2455, 3 => 3493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12157, 3 => 7405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6598, 3 => 11495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11805, 3 => 4455, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9625, 3 => 2090, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 4731, 3 => 2321, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 3578, 3 => 2608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 8504, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 4027, 3 => 1151, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5647, 3 => 4935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4219, 3 => 1870, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10968, 3 => 8054, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6970, 3 => 5447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3217, 3 => 5638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 8972, 3 => 669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5618, 3 => 12472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1457, 3 => 1280, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 8868, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8866, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 8371, 3 => 5972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 266, 3 => 4405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3706, 3 => 3244, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 6039, 3 => 5844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7200, 3 => 3283, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1502, 3 => 11282, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 12318, 3 => 2202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4523, 3 => 965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9587, 3 => 7011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2552, 3 => 2051, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12045, 3 => 10306, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 21, 2 => 11070, 3 => 5104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6627, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 23, 2 => 9889, 3 => 2121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 24, 2 => 829, 3 => 9701, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2201, 3 => 1819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6689, 3 => 12925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2139, 3 => 8757, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12004, 3 => 5948, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8704, 3 => 3191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8171, 3 => 10933, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6297, 3 => 7116, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 32, 2 => 616, 3 => 7146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 33, 2 => 5142, 3 => 9761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 34, 2 => 10377, 3 => 8138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7616, 3 => 5811, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7285, 3 => 9863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7764, 3 => 10867, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 12343, 3 => 9019, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4414, 3 => 8331, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3464, 3 => 642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6960, 3 => 2039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 786, 3 => 3021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 710, 3 => 2086, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 7423, 3 => 5601, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8120, 3 => 4885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 12385, 3 => 11990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9739, 3 => 10034, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 424, 3 => 10162, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1347, 3 => 7597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1450, 3 => 112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 7965, 3 => 8478, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8945, 3 => 7397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 6590, 3 => 8316, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6838, 3 => 9011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6174, 3 => 9410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 20, 2 => 255, 3 => 113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 21, 2 => 6197, 3 => 5835, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12902, 3 => 3844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 23, 2 => 4377, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 24, 2 => 5478, 3 => 8672, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4453, 3 => 2132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 26, 2 => 9724, 3 => 1380, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 27, 2 => 12131, 3 => 11526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12323, 3 => 9511, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8231, 3 => 1752, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 30, 2 => 497, 3 => 9022, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9288, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 32, 2 => 2481, 3 => 7515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 33, 2 => 2696, 3 => 268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 34, 2 => 4023, 3 => 12341, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7108, 3 => 5553, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C5_6.csv, table is 150x177 (3318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 5, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14, 13 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6 : integer_2d_array_t(0 to 149)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 4362, 3 => 416, 4 => 8909, 5 => 4156, 6 => 3216, 7 => 3112, 8 => 2560, 9 => 2912, 10 => 6405, 11 => 8593, 12 => 4969, 13 => 6723),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 2479, 3 => 1786, 4 => 8978, 5 => 3011, 6 => 4339, 7 => 9313, 8 => 6397, 9 => 2957, 10 => 7288, 11 => 5484, 12 => 6031, 13 => 10217),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 10175, 3 => 9009, 4 => 9889, 5 => 3091, 6 => 4985, 7 => 7267, 8 => 4092, 9 => 8874, 10 => 5671, 11 => 2777, 12 => 2189, 13 => 8716),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 9052, 3 => 4795, 4 => 3924, 5 => 3370, 6 => 10058, 7 => 1128, 8 => 9996, 9 => 10165, 10 => 9360, 11 => 4297, 12 => 434, 13 => 5138),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 2379, 3 => 7834, 4 => 4835, 5 => 2327, 6 => 9843, 7 => 804, 8 => 329, 9 => 8353, 10 => 7167, 11 => 3070, 12 => 1528, 13 => 7311),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 3435, 3 => 7871, 4 => 348, 5 => 3693, 6 => 1876, 7 => 6585, 8 => 10340, 9 => 7144, 10 => 5870, 11 => 2084, 12 => 4052, 13 => 2780),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 3917, 3 => 3111, 4 => 3476, 5 => 1304, 6 => 10331, 7 => 5939, 8 => 5199, 9 => 1611, 10 => 1991, 11 => 699, 12 => 8316, 13 => 9960),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 6883, 3 => 3237, 4 => 1717, 5 => 10752, 6 => 7891, 7 => 9764, 8 => 4745, 9 => 3888, 10 => 10009, 11 => 4176, 12 => 4614, 13 => 1567),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 10587, 3 => 2195, 4 => 1689, 5 => 2968, 6 => 5420, 7 => 2580, 8 => 2883, 9 => 6496, 10 => 111, 11 => 6023, 12 => 1024, 13 => 4449),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 3786, 3 => 8593, 4 => 2074, 5 => 3321, 6 => 5057, 7 => 1450, 8 => 3840, 9 => 5444, 10 => 6572, 11 => 3094, 12 => 9892, 13 => 1512),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 8548, 3 => 1848, 4 => 10372, 5 => 4585, 6 => 7313, 7 => 6536, 8 => 6379, 9 => 1766, 10 => 9462, 11 => 2456, 12 => 5606, 13 => 9975),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 8204, 3 => 10593, 4 => 7935, 5 => 3636, 6 => 3882, 7 => 394, 8 => 5968, 9 => 8561, 10 => 2395, 11 => 7289, 12 => 9267, 13 => 9978),
    12 => integer_vector_t'(0 => 13, 1 => 12, 2 => 7795, 3 => 74, 4 => 1633, 5 => 9542, 6 => 6867, 7 => 7352, 8 => 6417, 9 => 7568, 10 => 10623, 11 => 725, 12 => 2531, 13 => 9115),
    13 => integer_vector_t'(0 => 13, 1 => 13, 2 => 7151, 3 => 2482, 4 => 4260, 5 => 5003, 6 => 10105, 7 => 7419, 8 => 9203, 9 => 6691, 10 => 8798, 11 => 2092, 12 => 8263, 13 => 3755),
    14 => integer_vector_t'(0 => 13, 1 => 14, 2 => 3600, 3 => 570, 4 => 4527, 5 => 200, 6 => 9718, 7 => 6771, 8 => 1995, 9 => 8902, 10 => 5446, 11 => 768, 12 => 1103, 13 => 6520),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6304, 3 => 7621, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6498, 3 => 9209, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 7293, 3 => 6786, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5950, 3 => 1708, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8521, 3 => 1793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 6174, 3 => 7854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9773, 3 => 1190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9517, 3 => 10268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2181, 3 => 9349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 1949, 3 => 5560, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 1556, 3 => 555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8600, 3 => 3827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5072, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7928, 3 => 3542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3226, 3 => 3762, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7045, 3 => 2420, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9645, 3 => 2641, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2774, 3 => 2452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5331, 3 => 2031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9400, 3 => 7503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1850, 3 => 2338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10456, 3 => 9774, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1692, 3 => 9276, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 8, 2 => 10037, 3 => 4038, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3964, 3 => 338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 10, 2 => 2640, 3 => 5087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 11, 2 => 858, 3 => 3473, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5582, 3 => 5683, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9523, 3 => 916, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4107, 3 => 1559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4506, 3 => 3491, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8191, 3 => 4182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 17, 2 => 10192, 3 => 6157, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5668, 3 => 3305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3449, 3 => 1540, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4766, 3 => 2697, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4069, 3 => 6675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 22, 2 => 1117, 3 => 1016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5619, 3 => 3085, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8483, 3 => 8400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 25, 2 => 8255, 3 => 394, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6338, 3 => 5042, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 27, 2 => 6174, 3 => 5119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7203, 3 => 1989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 29, 2 => 1781, 3 => 5174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1464, 3 => 3559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3376, 3 => 4214, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7238, 3 => 67, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 10595, 3 => 8831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1221, 3 => 6513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5300, 3 => 4652, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1429, 3 => 9749, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7878, 3 => 5131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4435, 3 => 10284, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6331, 3 => 5507, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6662, 3 => 4941, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9614, 3 => 10238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 8400, 3 => 8025, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9156, 3 => 5630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7067, 3 => 8878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9027, 3 => 3415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1690, 3 => 3866, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2854, 3 => 8469, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6206, 3 => 630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 363, 3 => 5453, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4125, 3 => 7008, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1612, 3 => 6702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9069, 3 => 9226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5767, 3 => 4060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 3743, 3 => 9237, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7018, 3 => 5572, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8892, 3 => 4536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 853, 3 => 6064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8069, 3 => 5893, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2051, 3 => 2885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 10691, 3 => 3153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3602, 3 => 4055, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 328, 3 => 1717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2219, 3 => 9299, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1939, 3 => 7898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 617, 3 => 206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 8544, 3 => 1374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 10676, 3 => 3240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6672, 3 => 9489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3170, 3 => 7457, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7868, 3 => 5731, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6121, 3 => 10732, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4843, 3 => 9132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 580, 3 => 9591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 6267, 3 => 9290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3009, 3 => 2268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 195, 3 => 2419, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8016, 3 => 1557, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1516, 3 => 9195, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8062, 3 => 9064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 8968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 753, 3 => 7326, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6291, 3 => 3833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2614, 3 => 7844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2303, 3 => 646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2075, 3 => 611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4687, 3 => 362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 8684, 3 => 9940, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4830, 3 => 2065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7038, 3 => 1363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1769, 3 => 7837, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3801, 3 => 1689, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10070, 3 => 2359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3667, 3 => 9918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1914, 3 => 6920, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4244, 3 => 5669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10245, 3 => 7821, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7648, 3 => 3944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3310, 3 => 5488, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6346, 3 => 9666, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7088, 3 => 6122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1291, 3 => 7827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 10592, 3 => 8945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3609, 3 => 7120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 9168, 3 => 9112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6203, 3 => 8052, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3330, 3 => 2895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4264, 3 => 10563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10556, 3 => 6496, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8807, 3 => 7645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1999, 3 => 4530, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9202, 3 => 6818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3403, 3 => 1734, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2106, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 24, 2 => 6881, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 25, 2 => 3895, 3 => 2171, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4062, 3 => 6424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 27, 2 => 3755, 3 => 9536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4683, 3 => 2131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7347, 3 => 8027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C8_9.csv, table is 160x46 (920.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9 : integer_2d_array_t(0 to 159)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 6235, 3 => 2848, 4 => 3222),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5800, 3 => 3492, 4 => 5348),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2757, 3 => 927, 4 => 90),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6961, 3 => 4516, 4 => 4739),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1172, 3 => 3237, 4 => 6264),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1927, 3 => 2425, 4 => 3683),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3714, 3 => 6309, 4 => 2495),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 3070, 3 => 6342, 4 => 7154),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2428, 3 => 613, 4 => 3761),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 2906, 3 => 264, 4 => 5927),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 1716, 3 => 1950, 4 => 4273),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4613, 3 => 6179, 4 => 3491),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 4865, 3 => 3286, 4 => 6005),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1343, 3 => 5923, 4 => 3529),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 4589, 3 => 4035, 4 => 2132),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 1579, 3 => 3920, 4 => 6737),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1644, 3 => 1191, 4 => 5998),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 1482, 3 => 2381, 4 => 4620),
    18 => integer_vector_t'(0 => 4, 1 => 18, 2 => 6791, 3 => 6014, 4 => 6596),
    19 => integer_vector_t'(0 => 4, 1 => 19, 2 => 2738, 3 => 5918, 4 => 3786),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5156, 3 => 6166, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1504, 3 => 4356, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 130, 3 => 1904, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6027, 3 => 3187, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6718, 3 => 759, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6240, 3 => 2870, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2343, 3 => 1311, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1039, 3 => 5465, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6617, 3 => 2513, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1588, 3 => 5222, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6561, 3 => 535, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4765, 3 => 2054, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5966, 3 => 6892, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1969, 3 => 3869, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3571, 3 => 2420, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4632, 3 => 981, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3215, 3 => 4163, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 17, 2 => 973, 3 => 3117, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 18, 2 => 3802, 3 => 6198, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3794, 3 => 3948, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3196, 3 => 6126, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 1, 2 => 573, 3 => 1909, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 2, 2 => 850, 3 => 4034, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5622, 3 => 1601, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6005, 3 => 524, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5251, 3 => 5783, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 6, 2 => 172, 3 => 2032, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1875, 3 => 2475, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 8, 2 => 497, 3 => 1291, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2566, 3 => 3430, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1249, 3 => 740, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2944, 3 => 1948, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6528, 3 => 2899, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2243, 3 => 3616, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 14, 2 => 867, 3 => 3733, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1374, 3 => 4702, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4698, 3 => 2285, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4760, 3 => 3917, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1859, 3 => 4058, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6141, 3 => 3527, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2148, 3 => 5066, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1306, 3 => 145, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2319, 3 => 871, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3463, 3 => 1061, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5554, 3 => 6647, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5837, 3 => 339, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5821, 3 => 4932, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6356, 3 => 4756, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3930, 3 => 418, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 211, 3 => 3094, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1007, 3 => 4928, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3584, 3 => 1235, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6982, 3 => 2869, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1612, 3 => 1013, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 953, 3 => 4964, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4555, 3 => 4410, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4925, 3 => 4842, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5778, 3 => 600, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6509, 3 => 2417, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1260, 3 => 4903, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3369, 3 => 3031, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3557, 3 => 3224, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3028, 3 => 583, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3258, 3 => 440, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6226, 3 => 6655, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4895, 3 => 1094, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1481, 3 => 6847, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4433, 3 => 1932, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2107, 3 => 1649, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2119, 3 => 2065, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4003, 3 => 6388, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6720, 3 => 3622, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3694, 3 => 4521, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1164, 3 => 7050, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1965, 3 => 3613, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4331, 3 => 66, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2970, 3 => 1796, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4652, 3 => 3218, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1762, 3 => 4777, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5736, 3 => 1399, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 0, 2 => 970, 3 => 2572, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2062, 3 => 6599, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4597, 3 => 4870, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1228, 3 => 6913, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4159, 3 => 1037, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2916, 3 => 2362, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 6, 2 => 395, 3 => 1226, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6911, 3 => 4548, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4618, 3 => 2241, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4120, 3 => 4280, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5825, 3 => 474, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2154, 3 => 5558, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3793, 3 => 5471, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5707, 3 => 1595, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1403, 3 => 325, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6601, 3 => 5183, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6369, 3 => 4569, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4846, 3 => 896, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 18, 2 => 7092, 3 => 6184, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6764, 3 => 7127, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6358, 3 => 1951, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3117, 3 => 6960, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2710, 3 => 7062, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1133, 3 => 3604, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3694, 3 => 657, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1355, 3 => 110, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3329, 3 => 6736, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2505, 3 => 3407, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2462, 3 => 4806, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4216, 3 => 214, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5348, 3 => 5619, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6627, 3 => 6243, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 2644, 3 => 5073, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4212, 3 => 5088, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3463, 3 => 3889, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5306, 3 => 478, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4320, 3 => 6121, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3961, 3 => 1125, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5699, 3 => 1195, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6511, 3 => 792, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3934, 3 => 2778, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3238, 3 => 6587, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1111, 3 => 6596, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1457, 3 => 6226, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1446, 3 => 3885, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3907, 3 => 4043, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6839, 3 => 2873, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1733, 3 => 5615, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5202, 3 => 4269, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3024, 3 => 4722, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5445, 3 => 6372, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 11, 2 => 370, 3 => 1828, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4695, 3 => 1600, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 13, 2 => 680, 3 => 2074, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1801, 3 => 6690, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2669, 3 => 1377, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2463, 3 => 1681, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5972, 3 => 5171, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5728, 3 => 4284, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1696, 3 => 1459, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C9_10.csv, table is 162x46 (931.5 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10 : integer_2d_array_t(0 to 161)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 5611, 3 => 2563, 4 => 2900),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5220, 3 => 3143, 4 => 4813),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2481, 3 => 834, 4 => 81),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6265, 3 => 4064, 4 => 4265),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1055, 3 => 2914, 4 => 5638),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1734, 3 => 2182, 4 => 3315),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3342, 3 => 5678, 4 => 2246),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 2185, 3 => 552, 4 => 3385),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2615, 3 => 236, 4 => 5334),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 1546, 3 => 1755, 4 => 3846),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 4154, 3 => 5561, 4 => 3142),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4382, 3 => 2957, 4 => 5400),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 1209, 3 => 5329, 4 => 3179),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1421, 3 => 3528, 4 => 6063),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 1480, 3 => 1072, 4 => 5398),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 3843, 3 => 1777, 4 => 4369),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1334, 3 => 2145, 4 => 4163),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 2368, 3 => 5055, 4 => 260),
    18 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6118, 3 => 5405, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2994, 3 => 4370, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3405, 3 => 1669, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4640, 3 => 5550, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1354, 3 => 3921, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 5, 2 => 117, 3 => 1713, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5425, 3 => 2866, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6047, 3 => 683, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5616, 3 => 2582, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2108, 3 => 1179, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 10, 2 => 933, 3 => 4921, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5953, 3 => 2261, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1430, 3 => 4699, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5905, 3 => 480, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4289, 3 => 1846, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5374, 3 => 6208, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1775, 3 => 3476, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3216, 3 => 2178, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4165, 3 => 884, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2896, 3 => 3744, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 2801, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3423, 3 => 5579, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3404, 3 => 3552, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2876, 3 => 5515, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 516, 3 => 1719, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 765, 3 => 3631, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5059, 3 => 1441, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5629, 3 => 598, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5405, 3 => 473, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4724, 3 => 5210, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 155, 3 => 1832, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1689, 3 => 2229, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 449, 3 => 1164, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2308, 3 => 3088, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1122, 3 => 669, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2268, 3 => 5758, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5878, 3 => 2609, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 1, 2 => 782, 3 => 3359, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1231, 3 => 4231, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4225, 3 => 2052, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4286, 3 => 3517, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5531, 3 => 3184, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1935, 3 => 4560, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1174, 3 => 131, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3115, 3 => 956, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3129, 3 => 1088, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5238, 3 => 4440, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5722, 3 => 4280, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3540, 3 => 375, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 13, 2 => 191, 3 => 2782, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 14, 2 => 906, 3 => 4432, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3225, 3 => 1111, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6296, 3 => 2583, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1457, 3 => 903, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 855, 3 => 4475, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4097, 3 => 3970, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4433, 3 => 4361, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5198, 3 => 541, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1146, 3 => 4426, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3202, 3 => 2902, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2724, 3 => 525, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1083, 3 => 4124, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2326, 3 => 6003, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5605, 3 => 5990, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4376, 3 => 1579, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4407, 3 => 984, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1332, 3 => 6163, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5359, 3 => 3975, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1907, 3 => 1854, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3601, 3 => 5748, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6056, 3 => 3266, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3322, 3 => 4085, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1768, 3 => 3244, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2149, 3 => 144, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1589, 3 => 4291, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5154, 3 => 1252, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1855, 3 => 5939, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4820, 3 => 2706, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1475, 3 => 3360, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4266, 3 => 693, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4156, 3 => 2018, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2103, 3 => 752, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3710, 3 => 3853, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5123, 3 => 931, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6146, 3 => 3323, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1939, 3 => 5002, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5140, 3 => 1437, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1263, 3 => 293, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5949, 3 => 4665, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4548, 3 => 6380, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3171, 3 => 4690, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5204, 3 => 2114, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6384, 3 => 5565, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5722, 3 => 1757, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2805, 3 => 6264, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1202, 3 => 2616, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1018, 3 => 3244, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4018, 3 => 5289, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2257, 3 => 3067, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2483, 3 => 3073, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1196, 3 => 5329, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 649, 3 => 3918, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3791, 3 => 4581, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5028, 3 => 3803, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3119, 3 => 3506, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4779, 3 => 431, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3888, 3 => 5510, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4387, 3 => 4084, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5836, 3 => 1692, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5126, 3 => 1078, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 2, 2 => 5721, 3 => 6165, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3540, 3 => 2499, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2225, 3 => 6348, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1044, 3 => 1484, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6323, 3 => 4042, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1313, 3 => 5603, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1303, 3 => 3496, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3516, 3 => 3639, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5161, 3 => 2293, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4682, 3 => 3845, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3045, 3 => 643, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2818, 3 => 2616, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3267, 3 => 649, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6236, 3 => 593, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 16, 2 => 646, 3 => 2948, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4213, 3 => 1442, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5779, 3 => 1596, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2403, 3 => 1237, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2217, 3 => 1514, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5609, 3 => 716, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5155, 3 => 3858, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1517, 3 => 1312, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2554, 3 => 3158, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5280, 3 => 2643, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4990, 3 => 1353, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5648, 3 => 1170, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1152, 3 => 4366, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3561, 3 => 5368, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3581, 3 => 1411, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5647, 3 => 4661, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1542, 3 => 5401, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5078, 3 => 2687, 4 => -1),
    160 => integer_vector_t'(0 => 3, 1 => 16, 2 => 316, 3 => 1755, 4 => -1),
    161 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3392, 3 => 1991, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_2.csv, table is 20x100 (250.0 bytes)
  -- Resource estimation: 6 x 18 kB BRAMs or 3 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 5, 2 => 14, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_2 : integer_2d_array_t(0 to 19)(0 to 8) := (
    0 => integer_vector_t'(0 => 8, 1 => 20, 2 => 712, 3 => 2386, 4 => 6354, 5 => 4061, 6 => 1062, 7 => 5045, 8 => 5158),
    1 => integer_vector_t'(0 => 8, 1 => 21, 2 => 2543, 3 => 5748, 4 => 4822, 5 => 2348, 6 => 3089, 7 => 6328, 8 => 5876),
    2 => integer_vector_t'(0 => 8, 1 => 22, 2 => 926, 3 => 5701, 4 => 269, 5 => 3693, 6 => 2438, 7 => 3190, 8 => 3507),
    3 => integer_vector_t'(0 => 8, 1 => 23, 2 => 2802, 3 => 4520, 4 => 3577, 5 => 5324, 6 => 1091, 7 => 4667, 8 => 4449),
    4 => integer_vector_t'(0 => 8, 1 => 24, 2 => 5140, 3 => 2003, 4 => 1263, 5 => 4742, 6 => 6497, 7 => 1185, 8 => 6202),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4046, 3 => 6934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2855, 3 => 66, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6694, 3 => 212, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3439, 3 => 1158, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3850, 3 => 4422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5924, 3 => 290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1467, 3 => 4049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7820, 3 => 2242, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4606, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4633, 3 => 7877, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3884, 3 => 6868, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8935, 3 => 4996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3028, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5988, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7411, 3 => 3450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_3.csv, table is 15x170 (318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 13, 9 => 14, 10 => 14, 11 => 14, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_3 : integer_2d_array_t(0 to 14)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 416, 2 => 8909, 3 => 4156, 4 => 3216, 5 => 3112, 6 => 2560, 7 => 2912, 8 => 6405, 9 => 8593, 10 => 4969, 11 => 6723, 12 => 6912),
    1 => integer_vector_t'(0 => 12, 1 => 8978, 2 => 3011, 3 => 4339, 4 => 9312, 5 => 6396, 6 => 2957, 7 => 7288, 8 => 5485, 9 => 6031, 10 => 10218, 11 => 2226, 12 => 3575),
    2 => integer_vector_t'(0 => 12, 1 => 3383, 2 => 10059, 3 => 1114, 4 => 10008, 5 => 10147, 6 => 9384, 7 => 4290, 8 => 434, 9 => 5139, 10 => 3536, 11 => 1965, 12 => 2291),
    3 => integer_vector_t'(0 => 12, 1 => 2797, 2 => 3693, 3 => 7615, 4 => 7077, 5 => 743, 6 => 1941, 7 => 8716, 8 => 6215, 9 => 3840, 10 => 5140, 11 => 4582, 12 => 5420),
    4 => integer_vector_t'(0 => 12, 1 => 6110, 2 => 8551, 3 => 1515, 4 => 7404, 5 => 4879, 6 => 4946, 7 => 5383, 8 => 1831, 9 => 3441, 10 => 9569, 11 => 10472, 12 => 4306),
    5 => integer_vector_t'(0 => 3, 1 => 1505, 2 => 5682, 3 => 7778, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 7172, 2 => 6830, 3 => 6623, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7281, 2 => 3941, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 10270, 2 => 8669, 3 => 914, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 3622, 2 => 7563, 3 => 9388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 9930, 2 => 5058, 3 => 4554, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 4844, 2 => 9609, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 6883, 2 => 3237, 3 => 1714, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4768, 2 => 3878, 3 => 10017, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 10127, 2 => 3334, 3 => 8267, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_4.csv, table is 9x171 (192.375 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 13, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_4 : integer_2d_array_t(0 to 8)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 6295, 2 => 9626, 3 => 304, 4 => 7695, 5 => 4839, 6 => 4936, 7 => 1660, 8 => 144, 9 => 11203, 10 => 5567, 11 => 6347, 12 => 12557),
    1 => integer_vector_t'(0 => 12, 1 => 10691, 2 => 4988, 3 => 3859, 4 => 3734, 5 => 3071, 6 => 3494, 7 => 7687, 8 => 10313, 9 => 5964, 10 => 8069, 11 => 8296, 12 => 11090),
    2 => integer_vector_t'(0 => 12, 1 => 10774, 2 => 3613, 3 => 5208, 4 => 11177, 5 => 7676, 6 => 3549, 7 => 8746, 8 => 6583, 9 => 7239, 10 => 12265, 11 => 2674, 12 => 4292),
    3 => integer_vector_t'(0 => 12, 1 => 11869, 2 => 3708, 3 => 5981, 4 => 8718, 5 => 4908, 6 => 10650, 7 => 6805, 8 => 3334, 9 => 2627, 10 => 10461, 11 => 9285, 12 => 11120),
    4 => integer_vector_t'(0 => 3, 1 => 7844, 2 => 3079, 3 => 10773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 3385, 2 => 10854, 3 => 5747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1360, 2 => 12010, 3 => 12202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 6189, 2 => 4241, 3 => 2343, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9840, 2 => 12726, 3 => 4977, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_3.csv, table is 30x156 (585.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 13, 4 => 12, 5 => 12, 6 => 11, 7 => 12, 8 => 13, 9 => 12, 10 => 13, 11 => 12, 12 => 13, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_3 : integer_2d_array_t(0 to 29)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 2084, 3 => 1613, 4 => 1548, 5 => 1286, 6 => 1460, 7 => 3196, 8 => 4297, 9 => 2481, 10 => 3369, 11 => 3451, 12 => 4620, 13 => 2622),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 122, 3 => 1516, 4 => 3448, 5 => 2880, 6 => 1407, 7 => 1847, 8 => 3799, 9 => 3529, 10 => 373, 11 => 971, 12 => 4358, 13 => 3108),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 259, 3 => 3399, 4 => 929, 5 => 2650, 6 => 864, 7 => 3996, 8 => 3833, 9 => 107, 10 => 5287, 11 => 164, 12 => 3125, 13 => 2350),
    3 => integer_vector_t'(0 => 3, 1 => 3, 2 => 342, 3 => 3529, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4198, 3 => 2147, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1880, 3 => 4836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3864, 3 => 4910, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7, 2 => 243, 3 => 1542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3011, 3 => 1436, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2167, 3 => 2512, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4606, 3 => 1003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2835, 3 => 705, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3426, 3 => 2365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3848, 3 => 2474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1360, 3 => 1743, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 163, 3 => 2536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2583, 3 => 1180, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1542, 3 => 509, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4418, 3 => 1005, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5212, 3 => 5117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2155, 3 => 2922, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 347, 3 => 2696, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 226, 3 => 4296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1560, 3 => 487, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3926, 3 => 1640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 10, 2 => 149, 3 => 2928, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2364, 3 => 563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 12, 2 => 635, 3 => 688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 13, 2 => 231, 3 => 1684, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1129, 3 => 3894, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_5.csv, table is 18x168 (378.0 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 13, 8 => 13, 9 => 13, 10 => 14, 11 => 13, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_5 : integer_2d_array_t(0 to 17)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 5650, 2 => 4143, 3 => 8750, 4 => 583, 5 => 6720, 6 => 8071, 7 => 635, 8 => 1767, 9 => 1344, 10 => 6922, 11 => 738, 12 => 6658),
    1 => integer_vector_t'(0 => 12, 1 => 5696, 2 => 1685, 3 => 3207, 4 => 415, 5 => 7019, 6 => 5023, 7 => 5608, 8 => 2605, 9 => 857, 10 => 6915, 11 => 1770, 12 => 8016),
    2 => integer_vector_t'(0 => 12, 1 => 3992, 2 => 771, 3 => 2190, 4 => 7258, 5 => 8970, 6 => 7792, 7 => 1802, 8 => 1866, 9 => 6137, 10 => 8841, 11 => 886, 12 => 1931),
    3 => integer_vector_t'(0 => 12, 1 => 4108, 2 => 3781, 3 => 7577, 4 => 6810, 5 => 9322, 6 => 8226, 7 => 5396, 8 => 5867, 9 => 4428, 10 => 8827, 11 => 7766, 12 => 2254),
    4 => integer_vector_t'(0 => 12, 1 => 4247, 2 => 888, 3 => 4367, 4 => 8821, 5 => 9660, 6 => 324, 7 => 5864, 8 => 4774, 9 => 227, 10 => 7889, 11 => 6405, 12 => 8963),
    5 => integer_vector_t'(0 => 12, 1 => 9693, 2 => 500, 3 => 2520, 4 => 2227, 5 => 1811, 6 => 9330, 7 => 1928, 8 => 5140, 9 => 4030, 10 => 4824, 11 => 806, 12 => 3134),
    6 => integer_vector_t'(0 => 3, 1 => 1652, 2 => 8171, 3 => 1435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 3366, 2 => 6543, 3 => 3745, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9286, 2 => 8509, 3 => 4645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 7397, 2 => 5790, 3 => 8972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 6597, 2 => 4422, 3 => 1799, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 9276, 2 => 4041, 3 => 3847, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 8683, 2 => 7378, 3 => 4946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 5348, 2 => 1993, 3 => 9186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 6724, 2 => 9015, 3 => 5646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 4502, 2 => 4439, 3 => 8474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 5107, 2 => 7342, 3 => 9442, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 1387, 2 => 8910, 3 => 2660, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_4.csv, table is 33x133 (548.625 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 12, 4 => 13, 5 => 11, 6 => 10, 7 => 12, 8 => 11, 9 => 12, 10 => 10, 11 => 10, 12 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_4 : integer_2d_array_t(0 to 32)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 3, 2 => 3198, 3 => 478, 4 => 4207, 5 => 1481, 6 => 1009, 7 => 2616, 8 => 1924, 9 => 3437, 10 => 554, 11 => 683, 12 => 1801),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2681, 3 => 2135, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3107, 3 => 4027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2637, 3 => 3373, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 3830, 3 => 3449, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4129, 3 => 2060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4184, 3 => 2742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3946, 3 => 1070, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2239, 3 => 984, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1458, 3 => 3031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3003, 3 => 1328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1137, 3 => 1716, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 132, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1817, 3 => 638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1774, 3 => 3447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3632, 3 => 1257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 542, 3 => 3694, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1015, 3 => 1945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1948, 3 => 412, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 995, 3 => 2238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4141, 3 => 1907, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2480, 3 => 3079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3021, 3 => 1088, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 713, 3 => 1379, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 997, 3 => 3903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2323, 3 => 3361, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1110, 3 => 986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2532, 3 => 142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1690, 3 => 2405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1298, 3 => 1881, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 9, 2 => 615, 3 => 174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1648, 3 => 3112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1415, 3 => 2808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_5.csv, table is 27x160 (540.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 13, 2 => 13, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13, 9 => 13, 10 => 13, 11 => 13, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_5 : integer_2d_array_t(0 to 26)(0 to 12) := (
    0 => integer_vector_t'(0 => 12, 1 => 2765, 2 => 5713, 3 => 6426, 4 => 3596, 5 => 1374, 6 => 4811, 7 => 2182, 8 => 544, 9 => 3394, 10 => 2840, 11 => 4310, 12 => 771),
    1 => integer_vector_t'(0 => 12, 1 => 4951, 2 => 211, 3 => 2208, 4 => 723, 5 => 1246, 6 => 2928, 7 => 398, 8 => 5739, 9 => 265, 10 => 5601, 11 => 5993, 12 => 2615),
    2 => integer_vector_t'(0 => 12, 1 => 210, 2 => 4730, 3 => 5777, 4 => 3096, 5 => 4282, 6 => 6238, 7 => 4939, 8 => 1119, 9 => 6463, 10 => 5298, 11 => 6320, 12 => 4016),
    3 => integer_vector_t'(0 => 12, 1 => 4167, 2 => 2063, 3 => 4757, 4 => 3157, 5 => 5664, 6 => 3956, 7 => 6045, 8 => 563, 9 => 4284, 10 => 2441, 11 => 3412, 12 => 6334),
    4 => integer_vector_t'(0 => 12, 1 => 4201, 2 => 2428, 3 => 4474, 4 => 59, 5 => 1721, 6 => 736, 7 => 2997, 8 => 428, 9 => 3807, 10 => 1513, 11 => 4732, 12 => 6195),
    5 => integer_vector_t'(0 => 12, 1 => 2670, 2 => 3081, 3 => 5139, 4 => 3736, 5 => 1999, 6 => 5889, 7 => 4362, 8 => 3806, 9 => 4534, 10 => 5409, 11 => 6384, 12 => 5809),
    6 => integer_vector_t'(0 => 12, 1 => 5516, 2 => 1622, 3 => 2906, 4 => 3285, 5 => 1257, 6 => 5797, 7 => 3816, 8 => 817, 9 => 875, 10 => 2311, 11 => 3543, 12 => 1205),
    7 => integer_vector_t'(0 => 12, 1 => 4244, 2 => 2184, 3 => 5415, 4 => 1705, 5 => 5642, 6 => 4886, 7 => 2333, 8 => 287, 9 => 1848, 10 => 1121, 11 => 3595, 12 => 6022),
    8 => integer_vector_t'(0 => 12, 1 => 2142, 2 => 2830, 3 => 4069, 4 => 5654, 5 => 1295, 6 => 2951, 7 => 3919, 8 => 1356, 9 => 884, 10 => 1786, 11 => 396, 12 => 4738),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2161, 3 => 2653, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1380, 3 => 1461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2502, 3 => 3707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3971, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5985, 3 => 6062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1733, 3 => 6028, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3786, 3 => 1936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4292, 3 => 956, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5692, 3 => 3417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 266, 3 => 4878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4913, 3 => 3247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4763, 3 => 3937, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3590, 3 => 2903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2566, 3 => 4215, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5208, 3 => 4707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3940, 3 => 3388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5109, 3 => 4556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4908, 3 => 4177, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C4_5.csv, table is 35x30 (131.25 bytes)
  -- Resource estimation: 2 x 18 kB BRAMs or 1 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 4, 2 => 12, 3 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C4_5 : integer_2d_array_t(0 to 34)(0 to 3) := (
    0 => integer_vector_t'(0 => 3, 1 => 5, 2 => 896, 3 => 1565),
    1 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2493, 3 => 184),
    2 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 3210),
    3 => integer_vector_t'(0 => 3, 1 => 8, 2 => 727, 3 => 1339),
    4 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3428, 3 => 612),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2663, 3 => 1947),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 230, 3 => 2695),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2025, 3 => 2794),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3039, 3 => 283),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 862, 3 => 2889),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 376, 3 => 2110),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2034, 3 => 2286),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 951, 3 => 2068),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3108, 3 => 3542),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 307, 3 => 1421),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2272, 3 => 1197),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1800, 3 => 3280),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 331, 3 => 2308),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 465, 3 => 2552),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1038, 3 => 2479),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1383, 3 => 343),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 94, 3 => 236),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2619, 3 => 121),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1497, 3 => 2774),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2116, 3 => 1855),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 722, 3 => 1584),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2767, 3 => 1881),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2701, 3 => 1610),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3283, 3 => 1732),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 168, 3 => 1099),
    30 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3074, 3 => 243),
    31 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3460, 3 => 945),
    32 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2049, 3 => 1746),
    33 => integer_vector_t'(0 => 3, 1 => 8, 2 => 566, 3 => 1427),
    34 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3545, 3 => 1168)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C5_6.csv, table is 37x139 (642.875 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 3, 2 => 12, 3 => 12, 4 => 11, 5 => 10, 6 => 10, 7 => 10, 8 => 11, 9 => 9, 10 => 12, 11 => 12, 12 => 11, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C5_6 : integer_2d_array_t(0 to 36)(0 to 13) := (
    0 => integer_vector_t'(0 => 13, 1 => 3, 2 => 2409, 3 => 499, 4 => 1481, 5 => 908, 6 => 559, 7 => 716, 8 => 1270, 9 => 333, 10 => 2508, 11 => 2264, 12 => 1702, 13 => 2805),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2447, 3 => 1926, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 414, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2114, 3 => 842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 573, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2383, 3 => 2112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2286, 3 => 2348, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 545, 3 => 819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1264, 3 => 143, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1701, 3 => 2258, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 964, 3 => 166, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 114, 3 => 2413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2243, 3 => 81, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1245, 3 => 1581, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 1, 2 => 775, 3 => 169, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1696, 3 => 1104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1914, 3 => 2831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 4, 2 => 532, 3 => 1450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 5, 2 => 91, 3 => 974, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 6, 2 => 497, 3 => 2228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2326, 3 => 1579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2482, 3 => 256, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1117, 3 => 1261, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1257, 3 => 1658, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1478, 3 => 1225, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2511, 3 => 980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2320, 3 => 2675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 435, 3 => 1278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 228, 3 => 503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1885, 3 => 2369, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 1, 2 => 57, 3 => 483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 2, 2 => 838, 3 => 1050, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1231, 3 => 1990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1738, 3 => 68, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2392, 3 => 951, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 6, 2 => 163, 3 => 645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2644, 3 => 1704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C8_9.csv, table is 40x37 (185.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 2, 2 => 11, 3 => 11, 4 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C8_9 : integer_2d_array_t(0 to 39)(0 to 4) := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 1558, 3 => 712, 4 => 805),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 1450, 3 => 873, 4 => 1337),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 1741, 3 => 1129, 4 => 1184),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 294, 3 => 806, 4 => 1566),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 482, 3 => 605, 4 => 923),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 926, 3 => 1578, 4 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 777, 3 => 1374, 4 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 608, 3 => 151, 4 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1195, 3 => 210, 4 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1484, 3 => 692, 4 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 0, 2 => 427, 3 => 488, 4 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 1, 2 => 828, 3 => 1124, 4 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 1366, 4 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1500, 3 => 835, 4 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1496, 3 => 502, 4 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1006, 3 => 1701, 4 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1155, 3 => 97, 4 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 657, 3 => 1403, 4 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1453, 3 => 624, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 429, 3 => 1495, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 809, 3 => 385, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 367, 3 => 151, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1323, 3 => 202, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 960, 3 => 318, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1451, 3 => 1039, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1098, 3 => 1722, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1015, 3 => 1428, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1261, 3 => 1564, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 544, 3 => 1190, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1472, 3 => 1246, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 508, 3 => 630, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 421, 3 => 1704, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 284, 3 => 898, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 392, 3 => 577, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1155, 3 => 556, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 0, 2 => 631, 3 => 1000, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 1, 2 => 732, 3 => 1368, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1328, 3 => 329, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1515, 3 => 506, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1104, 3 => 1172, 4 => -1)
  );


  -- Record with LDPC metadata
  type ldpc_metadata_t is record
    addr : integer;
    q : integer;
    stage_0_loops: integer;
    stage_0_rows: integer;
    stage_1_loops: integer;
    stage_1_rows: integer;
  end record ldpc_metadata_t;

  -- Reduce the footprint of this
  constant LDPC_TABLE_DATA_WIDTH : integer := numbits(max(DVB_N_LDPC));

  -- Use this function to get the starting address of a given config within the LDPC_DATA_TABLE
  function get_ldpc_metadata (
    constant frame_length : frame_type_t;
    constant code_rate : code_rate_t) return ldpc_metadata_t;


  constant LDPC_DATA_TABLE : std_logic_vector_2d_t(0 to 6446)(LDPC_TABLE_DATA_WIDTH - 1 downto 0) := (
    -- Table for fecframe_normal, C1_2
    0 => std_logic_vector(to_unsigned(54, LDPC_TABLE_DATA_WIDTH)),
    1 => std_logic_vector(to_unsigned(9318, LDPC_TABLE_DATA_WIDTH)),
    2 => std_logic_vector(to_unsigned(14392, LDPC_TABLE_DATA_WIDTH)),
    3 => std_logic_vector(to_unsigned(27561, LDPC_TABLE_DATA_WIDTH)),
    4 => std_logic_vector(to_unsigned(26909, LDPC_TABLE_DATA_WIDTH)),
    5 => std_logic_vector(to_unsigned(10219, LDPC_TABLE_DATA_WIDTH)),
    6 => std_logic_vector(to_unsigned(2534, LDPC_TABLE_DATA_WIDTH)),
    7 => std_logic_vector(to_unsigned(8597, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    8 => std_logic_vector(to_unsigned(55, LDPC_TABLE_DATA_WIDTH)),
    9 => std_logic_vector(to_unsigned(7263, LDPC_TABLE_DATA_WIDTH)),
    10 => std_logic_vector(to_unsigned(4635, LDPC_TABLE_DATA_WIDTH)),
    11 => std_logic_vector(to_unsigned(2530, LDPC_TABLE_DATA_WIDTH)),
    12 => std_logic_vector(to_unsigned(28130, LDPC_TABLE_DATA_WIDTH)),
    13 => std_logic_vector(to_unsigned(3033, LDPC_TABLE_DATA_WIDTH)),
    14 => std_logic_vector(to_unsigned(23830, LDPC_TABLE_DATA_WIDTH)),
    15 => std_logic_vector(to_unsigned(3651, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    16 => std_logic_vector(to_unsigned(56, LDPC_TABLE_DATA_WIDTH)),
    17 => std_logic_vector(to_unsigned(24731, LDPC_TABLE_DATA_WIDTH)),
    18 => std_logic_vector(to_unsigned(23583, LDPC_TABLE_DATA_WIDTH)),
    19 => std_logic_vector(to_unsigned(26036, LDPC_TABLE_DATA_WIDTH)),
    20 => std_logic_vector(to_unsigned(17299, LDPC_TABLE_DATA_WIDTH)),
    21 => std_logic_vector(to_unsigned(5750, LDPC_TABLE_DATA_WIDTH)),
    22 => std_logic_vector(to_unsigned(792, LDPC_TABLE_DATA_WIDTH)),
    23 => std_logic_vector(to_unsigned(9169, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    24 => std_logic_vector(to_unsigned(57, LDPC_TABLE_DATA_WIDTH)),
    25 => std_logic_vector(to_unsigned(5811, LDPC_TABLE_DATA_WIDTH)),
    26 => std_logic_vector(to_unsigned(26154, LDPC_TABLE_DATA_WIDTH)),
    27 => std_logic_vector(to_unsigned(18653, LDPC_TABLE_DATA_WIDTH)),
    28 => std_logic_vector(to_unsigned(11551, LDPC_TABLE_DATA_WIDTH)),
    29 => std_logic_vector(to_unsigned(15447, LDPC_TABLE_DATA_WIDTH)),
    30 => std_logic_vector(to_unsigned(13685, LDPC_TABLE_DATA_WIDTH)),
    31 => std_logic_vector(to_unsigned(16264, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    32 => std_logic_vector(to_unsigned(58, LDPC_TABLE_DATA_WIDTH)),
    33 => std_logic_vector(to_unsigned(12610, LDPC_TABLE_DATA_WIDTH)),
    34 => std_logic_vector(to_unsigned(11347, LDPC_TABLE_DATA_WIDTH)),
    35 => std_logic_vector(to_unsigned(28768, LDPC_TABLE_DATA_WIDTH)),
    36 => std_logic_vector(to_unsigned(2792, LDPC_TABLE_DATA_WIDTH)),
    37 => std_logic_vector(to_unsigned(3174, LDPC_TABLE_DATA_WIDTH)),
    38 => std_logic_vector(to_unsigned(29371, LDPC_TABLE_DATA_WIDTH)),
    39 => std_logic_vector(to_unsigned(12997, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    40 => std_logic_vector(to_unsigned(59, LDPC_TABLE_DATA_WIDTH)),
    41 => std_logic_vector(to_unsigned(16789, LDPC_TABLE_DATA_WIDTH)),
    42 => std_logic_vector(to_unsigned(16018, LDPC_TABLE_DATA_WIDTH)),
    43 => std_logic_vector(to_unsigned(21449, LDPC_TABLE_DATA_WIDTH)),
    44 => std_logic_vector(to_unsigned(6165, LDPC_TABLE_DATA_WIDTH)),
    45 => std_logic_vector(to_unsigned(21202, LDPC_TABLE_DATA_WIDTH)),
    46 => std_logic_vector(to_unsigned(15850, LDPC_TABLE_DATA_WIDTH)),
    47 => std_logic_vector(to_unsigned(3186, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    48 => std_logic_vector(to_unsigned(60, LDPC_TABLE_DATA_WIDTH)),
    49 => std_logic_vector(to_unsigned(31016, LDPC_TABLE_DATA_WIDTH)),
    50 => std_logic_vector(to_unsigned(21449, LDPC_TABLE_DATA_WIDTH)),
    51 => std_logic_vector(to_unsigned(17618, LDPC_TABLE_DATA_WIDTH)),
    52 => std_logic_vector(to_unsigned(6213, LDPC_TABLE_DATA_WIDTH)),
    53 => std_logic_vector(to_unsigned(12166, LDPC_TABLE_DATA_WIDTH)),
    54 => std_logic_vector(to_unsigned(8334, LDPC_TABLE_DATA_WIDTH)),
    55 => std_logic_vector(to_unsigned(18212, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    56 => std_logic_vector(to_unsigned(61, LDPC_TABLE_DATA_WIDTH)),
    57 => std_logic_vector(to_unsigned(22836, LDPC_TABLE_DATA_WIDTH)),
    58 => std_logic_vector(to_unsigned(14213, LDPC_TABLE_DATA_WIDTH)),
    59 => std_logic_vector(to_unsigned(11327, LDPC_TABLE_DATA_WIDTH)),
    60 => std_logic_vector(to_unsigned(5896, LDPC_TABLE_DATA_WIDTH)),
    61 => std_logic_vector(to_unsigned(718, LDPC_TABLE_DATA_WIDTH)),
    62 => std_logic_vector(to_unsigned(11727, LDPC_TABLE_DATA_WIDTH)),
    63 => std_logic_vector(to_unsigned(9308, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    64 => std_logic_vector(to_unsigned(62, LDPC_TABLE_DATA_WIDTH)),
    65 => std_logic_vector(to_unsigned(2091, LDPC_TABLE_DATA_WIDTH)),
    66 => std_logic_vector(to_unsigned(24941, LDPC_TABLE_DATA_WIDTH)),
    67 => std_logic_vector(to_unsigned(29966, LDPC_TABLE_DATA_WIDTH)),
    68 => std_logic_vector(to_unsigned(23634, LDPC_TABLE_DATA_WIDTH)),
    69 => std_logic_vector(to_unsigned(9013, LDPC_TABLE_DATA_WIDTH)),
    70 => std_logic_vector(to_unsigned(15587, LDPC_TABLE_DATA_WIDTH)),
    71 => std_logic_vector(to_unsigned(5444, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    72 => std_logic_vector(to_unsigned(63, LDPC_TABLE_DATA_WIDTH)),
    73 => std_logic_vector(to_unsigned(22207, LDPC_TABLE_DATA_WIDTH)),
    74 => std_logic_vector(to_unsigned(3983, LDPC_TABLE_DATA_WIDTH)),
    75 => std_logic_vector(to_unsigned(16904, LDPC_TABLE_DATA_WIDTH)),
    76 => std_logic_vector(to_unsigned(28534, LDPC_TABLE_DATA_WIDTH)),
    77 => std_logic_vector(to_unsigned(21415, LDPC_TABLE_DATA_WIDTH)),
    78 => std_logic_vector(to_unsigned(27524, LDPC_TABLE_DATA_WIDTH)),
    79 => std_logic_vector(to_unsigned(25912, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    80 => std_logic_vector(to_unsigned(64, LDPC_TABLE_DATA_WIDTH)),
    81 => std_logic_vector(to_unsigned(25687, LDPC_TABLE_DATA_WIDTH)),
    82 => std_logic_vector(to_unsigned(4501, LDPC_TABLE_DATA_WIDTH)),
    83 => std_logic_vector(to_unsigned(22193, LDPC_TABLE_DATA_WIDTH)),
    84 => std_logic_vector(to_unsigned(14665, LDPC_TABLE_DATA_WIDTH)),
    85 => std_logic_vector(to_unsigned(14798, LDPC_TABLE_DATA_WIDTH)),
    86 => std_logic_vector(to_unsigned(16158, LDPC_TABLE_DATA_WIDTH)),
    87 => std_logic_vector(to_unsigned(5491, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    88 => std_logic_vector(to_unsigned(65, LDPC_TABLE_DATA_WIDTH)),
    89 => std_logic_vector(to_unsigned(4520, LDPC_TABLE_DATA_WIDTH)),
    90 => std_logic_vector(to_unsigned(17094, LDPC_TABLE_DATA_WIDTH)),
    91 => std_logic_vector(to_unsigned(23397, LDPC_TABLE_DATA_WIDTH)),
    92 => std_logic_vector(to_unsigned(4264, LDPC_TABLE_DATA_WIDTH)),
    93 => std_logic_vector(to_unsigned(22370, LDPC_TABLE_DATA_WIDTH)),
    94 => std_logic_vector(to_unsigned(16941, LDPC_TABLE_DATA_WIDTH)),
    95 => std_logic_vector(to_unsigned(21526, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    96 => std_logic_vector(to_unsigned(66, LDPC_TABLE_DATA_WIDTH)),
    97 => std_logic_vector(to_unsigned(10490, LDPC_TABLE_DATA_WIDTH)),
    98 => std_logic_vector(to_unsigned(6182, LDPC_TABLE_DATA_WIDTH)),
    99 => std_logic_vector(to_unsigned(32370, LDPC_TABLE_DATA_WIDTH)),
    100 => std_logic_vector(to_unsigned(9597, LDPC_TABLE_DATA_WIDTH)),
    101 => std_logic_vector(to_unsigned(30841, LDPC_TABLE_DATA_WIDTH)),
    102 => std_logic_vector(to_unsigned(25954, LDPC_TABLE_DATA_WIDTH)),
    103 => std_logic_vector(to_unsigned(2762, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    104 => std_logic_vector(to_unsigned(67, LDPC_TABLE_DATA_WIDTH)),
    105 => std_logic_vector(to_unsigned(22120, LDPC_TABLE_DATA_WIDTH)),
    106 => std_logic_vector(to_unsigned(22865, LDPC_TABLE_DATA_WIDTH)),
    107 => std_logic_vector(to_unsigned(29870, LDPC_TABLE_DATA_WIDTH)),
    108 => std_logic_vector(to_unsigned(15147, LDPC_TABLE_DATA_WIDTH)),
    109 => std_logic_vector(to_unsigned(13668, LDPC_TABLE_DATA_WIDTH)),
    110 => std_logic_vector(to_unsigned(14955, LDPC_TABLE_DATA_WIDTH)),
    111 => std_logic_vector(to_unsigned(19235, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    112 => std_logic_vector(to_unsigned(68, LDPC_TABLE_DATA_WIDTH)),
    113 => std_logic_vector(to_unsigned(6689, LDPC_TABLE_DATA_WIDTH)),
    114 => std_logic_vector(to_unsigned(18408, LDPC_TABLE_DATA_WIDTH)),
    115 => std_logic_vector(to_unsigned(18346, LDPC_TABLE_DATA_WIDTH)),
    116 => std_logic_vector(to_unsigned(9918, LDPC_TABLE_DATA_WIDTH)),
    117 => std_logic_vector(to_unsigned(25746, LDPC_TABLE_DATA_WIDTH)),
    118 => std_logic_vector(to_unsigned(5443, LDPC_TABLE_DATA_WIDTH)),
    119 => std_logic_vector(to_unsigned(20645, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    120 => std_logic_vector(to_unsigned(69, LDPC_TABLE_DATA_WIDTH)),
    121 => std_logic_vector(to_unsigned(29982, LDPC_TABLE_DATA_WIDTH)),
    122 => std_logic_vector(to_unsigned(12529, LDPC_TABLE_DATA_WIDTH)),
    123 => std_logic_vector(to_unsigned(13858, LDPC_TABLE_DATA_WIDTH)),
    124 => std_logic_vector(to_unsigned(4746, LDPC_TABLE_DATA_WIDTH)),
    125 => std_logic_vector(to_unsigned(30370, LDPC_TABLE_DATA_WIDTH)),
    126 => std_logic_vector(to_unsigned(10023, LDPC_TABLE_DATA_WIDTH)),
    127 => std_logic_vector(to_unsigned(24828, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    128 => std_logic_vector(to_unsigned(70, LDPC_TABLE_DATA_WIDTH)),
    129 => std_logic_vector(to_unsigned(1262, LDPC_TABLE_DATA_WIDTH)),
    130 => std_logic_vector(to_unsigned(28032, LDPC_TABLE_DATA_WIDTH)),
    131 => std_logic_vector(to_unsigned(29888, LDPC_TABLE_DATA_WIDTH)),
    132 => std_logic_vector(to_unsigned(13063, LDPC_TABLE_DATA_WIDTH)),
    133 => std_logic_vector(to_unsigned(24033, LDPC_TABLE_DATA_WIDTH)),
    134 => std_logic_vector(to_unsigned(21951, LDPC_TABLE_DATA_WIDTH)),
    135 => std_logic_vector(to_unsigned(7863, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    136 => std_logic_vector(to_unsigned(71, LDPC_TABLE_DATA_WIDTH)),
    137 => std_logic_vector(to_unsigned(6594, LDPC_TABLE_DATA_WIDTH)),
    138 => std_logic_vector(to_unsigned(29642, LDPC_TABLE_DATA_WIDTH)),
    139 => std_logic_vector(to_unsigned(31451, LDPC_TABLE_DATA_WIDTH)),
    140 => std_logic_vector(to_unsigned(14831, LDPC_TABLE_DATA_WIDTH)),
    141 => std_logic_vector(to_unsigned(9509, LDPC_TABLE_DATA_WIDTH)),
    142 => std_logic_vector(to_unsigned(9335, LDPC_TABLE_DATA_WIDTH)),
    143 => std_logic_vector(to_unsigned(31552, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    144 => std_logic_vector(to_unsigned(72, LDPC_TABLE_DATA_WIDTH)),
    145 => std_logic_vector(to_unsigned(1358, LDPC_TABLE_DATA_WIDTH)),
    146 => std_logic_vector(to_unsigned(6454, LDPC_TABLE_DATA_WIDTH)),
    147 => std_logic_vector(to_unsigned(16633, LDPC_TABLE_DATA_WIDTH)),
    148 => std_logic_vector(to_unsigned(20354, LDPC_TABLE_DATA_WIDTH)),
    149 => std_logic_vector(to_unsigned(24598, LDPC_TABLE_DATA_WIDTH)),
    150 => std_logic_vector(to_unsigned(624, LDPC_TABLE_DATA_WIDTH)),
    151 => std_logic_vector(to_unsigned(5265, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    152 => std_logic_vector(to_unsigned(73, LDPC_TABLE_DATA_WIDTH)),
    153 => std_logic_vector(to_unsigned(19529, LDPC_TABLE_DATA_WIDTH)),
    154 => std_logic_vector(to_unsigned(295, LDPC_TABLE_DATA_WIDTH)),
    155 => std_logic_vector(to_unsigned(18011, LDPC_TABLE_DATA_WIDTH)),
    156 => std_logic_vector(to_unsigned(3080, LDPC_TABLE_DATA_WIDTH)),
    157 => std_logic_vector(to_unsigned(13364, LDPC_TABLE_DATA_WIDTH)),
    158 => std_logic_vector(to_unsigned(8032, LDPC_TABLE_DATA_WIDTH)),
    159 => std_logic_vector(to_unsigned(15323, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    160 => std_logic_vector(to_unsigned(74, LDPC_TABLE_DATA_WIDTH)),
    161 => std_logic_vector(to_unsigned(11981, LDPC_TABLE_DATA_WIDTH)),
    162 => std_logic_vector(to_unsigned(1510, LDPC_TABLE_DATA_WIDTH)),
    163 => std_logic_vector(to_unsigned(7960, LDPC_TABLE_DATA_WIDTH)),
    164 => std_logic_vector(to_unsigned(21462, LDPC_TABLE_DATA_WIDTH)),
    165 => std_logic_vector(to_unsigned(9129, LDPC_TABLE_DATA_WIDTH)),
    166 => std_logic_vector(to_unsigned(11370, LDPC_TABLE_DATA_WIDTH)),
    167 => std_logic_vector(to_unsigned(25741, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    168 => std_logic_vector(to_unsigned(75, LDPC_TABLE_DATA_WIDTH)),
    169 => std_logic_vector(to_unsigned(9276, LDPC_TABLE_DATA_WIDTH)),
    170 => std_logic_vector(to_unsigned(29656, LDPC_TABLE_DATA_WIDTH)),
    171 => std_logic_vector(to_unsigned(4543, LDPC_TABLE_DATA_WIDTH)),
    172 => std_logic_vector(to_unsigned(30699, LDPC_TABLE_DATA_WIDTH)),
    173 => std_logic_vector(to_unsigned(20646, LDPC_TABLE_DATA_WIDTH)),
    174 => std_logic_vector(to_unsigned(21921, LDPC_TABLE_DATA_WIDTH)),
    175 => std_logic_vector(to_unsigned(28050, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    176 => std_logic_vector(to_unsigned(76, LDPC_TABLE_DATA_WIDTH)),
    177 => std_logic_vector(to_unsigned(15975, LDPC_TABLE_DATA_WIDTH)),
    178 => std_logic_vector(to_unsigned(25634, LDPC_TABLE_DATA_WIDTH)),
    179 => std_logic_vector(to_unsigned(5520, LDPC_TABLE_DATA_WIDTH)),
    180 => std_logic_vector(to_unsigned(31119, LDPC_TABLE_DATA_WIDTH)),
    181 => std_logic_vector(to_unsigned(13715, LDPC_TABLE_DATA_WIDTH)),
    182 => std_logic_vector(to_unsigned(21949, LDPC_TABLE_DATA_WIDTH)),
    183 => std_logic_vector(to_unsigned(19605, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    184 => std_logic_vector(to_unsigned(77, LDPC_TABLE_DATA_WIDTH)),
    185 => std_logic_vector(to_unsigned(18688, LDPC_TABLE_DATA_WIDTH)),
    186 => std_logic_vector(to_unsigned(4608, LDPC_TABLE_DATA_WIDTH)),
    187 => std_logic_vector(to_unsigned(31755, LDPC_TABLE_DATA_WIDTH)),
    188 => std_logic_vector(to_unsigned(30165, LDPC_TABLE_DATA_WIDTH)),
    189 => std_logic_vector(to_unsigned(13103, LDPC_TABLE_DATA_WIDTH)),
    190 => std_logic_vector(to_unsigned(10706, LDPC_TABLE_DATA_WIDTH)),
    191 => std_logic_vector(to_unsigned(29224, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    192 => std_logic_vector(to_unsigned(78, LDPC_TABLE_DATA_WIDTH)),
    193 => std_logic_vector(to_unsigned(21514, LDPC_TABLE_DATA_WIDTH)),
    194 => std_logic_vector(to_unsigned(23117, LDPC_TABLE_DATA_WIDTH)),
    195 => std_logic_vector(to_unsigned(12245, LDPC_TABLE_DATA_WIDTH)),
    196 => std_logic_vector(to_unsigned(26035, LDPC_TABLE_DATA_WIDTH)),
    197 => std_logic_vector(to_unsigned(31656, LDPC_TABLE_DATA_WIDTH)),
    198 => std_logic_vector(to_unsigned(25631, LDPC_TABLE_DATA_WIDTH)),
    199 => std_logic_vector(to_unsigned(30699, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    200 => std_logic_vector(to_unsigned(79, LDPC_TABLE_DATA_WIDTH)),
    201 => std_logic_vector(to_unsigned(9674, LDPC_TABLE_DATA_WIDTH)),
    202 => std_logic_vector(to_unsigned(24966, LDPC_TABLE_DATA_WIDTH)),
    203 => std_logic_vector(to_unsigned(31285, LDPC_TABLE_DATA_WIDTH)),
    204 => std_logic_vector(to_unsigned(29908, LDPC_TABLE_DATA_WIDTH)),
    205 => std_logic_vector(to_unsigned(17042, LDPC_TABLE_DATA_WIDTH)),
    206 => std_logic_vector(to_unsigned(24588, LDPC_TABLE_DATA_WIDTH)),
    207 => std_logic_vector(to_unsigned(31857, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    208 => std_logic_vector(to_unsigned(80, LDPC_TABLE_DATA_WIDTH)),
    209 => std_logic_vector(to_unsigned(21856, LDPC_TABLE_DATA_WIDTH)),
    210 => std_logic_vector(to_unsigned(27777, LDPC_TABLE_DATA_WIDTH)),
    211 => std_logic_vector(to_unsigned(29919, LDPC_TABLE_DATA_WIDTH)),
    212 => std_logic_vector(to_unsigned(27000, LDPC_TABLE_DATA_WIDTH)),
    213 => std_logic_vector(to_unsigned(14897, LDPC_TABLE_DATA_WIDTH)),
    214 => std_logic_vector(to_unsigned(11409, LDPC_TABLE_DATA_WIDTH)),
    215 => std_logic_vector(to_unsigned(7122, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    216 => std_logic_vector(to_unsigned(81, LDPC_TABLE_DATA_WIDTH)),
    217 => std_logic_vector(to_unsigned(29773, LDPC_TABLE_DATA_WIDTH)),
    218 => std_logic_vector(to_unsigned(23310, LDPC_TABLE_DATA_WIDTH)),
    219 => std_logic_vector(to_unsigned(263, LDPC_TABLE_DATA_WIDTH)),
    220 => std_logic_vector(to_unsigned(4877, LDPC_TABLE_DATA_WIDTH)),
    221 => std_logic_vector(to_unsigned(28622, LDPC_TABLE_DATA_WIDTH)),
    222 => std_logic_vector(to_unsigned(20545, LDPC_TABLE_DATA_WIDTH)),
    223 => std_logic_vector(to_unsigned(22092, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    224 => std_logic_vector(to_unsigned(82, LDPC_TABLE_DATA_WIDTH)),
    225 => std_logic_vector(to_unsigned(15605, LDPC_TABLE_DATA_WIDTH)),
    226 => std_logic_vector(to_unsigned(5651, LDPC_TABLE_DATA_WIDTH)),
    227 => std_logic_vector(to_unsigned(21864, LDPC_TABLE_DATA_WIDTH)),
    228 => std_logic_vector(to_unsigned(3967, LDPC_TABLE_DATA_WIDTH)),
    229 => std_logic_vector(to_unsigned(14419, LDPC_TABLE_DATA_WIDTH)),
    230 => std_logic_vector(to_unsigned(22757, LDPC_TABLE_DATA_WIDTH)),
    231 => std_logic_vector(to_unsigned(15896, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    232 => std_logic_vector(to_unsigned(83, LDPC_TABLE_DATA_WIDTH)),
    233 => std_logic_vector(to_unsigned(30145, LDPC_TABLE_DATA_WIDTH)),
    234 => std_logic_vector(to_unsigned(1759, LDPC_TABLE_DATA_WIDTH)),
    235 => std_logic_vector(to_unsigned(10139, LDPC_TABLE_DATA_WIDTH)),
    236 => std_logic_vector(to_unsigned(29223, LDPC_TABLE_DATA_WIDTH)),
    237 => std_logic_vector(to_unsigned(26086, LDPC_TABLE_DATA_WIDTH)),
    238 => std_logic_vector(to_unsigned(10556, LDPC_TABLE_DATA_WIDTH)),
    239 => std_logic_vector(to_unsigned(5098, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    240 => std_logic_vector(to_unsigned(84, LDPC_TABLE_DATA_WIDTH)),
    241 => std_logic_vector(to_unsigned(18815, LDPC_TABLE_DATA_WIDTH)),
    242 => std_logic_vector(to_unsigned(16575, LDPC_TABLE_DATA_WIDTH)),
    243 => std_logic_vector(to_unsigned(2936, LDPC_TABLE_DATA_WIDTH)),
    244 => std_logic_vector(to_unsigned(24457, LDPC_TABLE_DATA_WIDTH)),
    245 => std_logic_vector(to_unsigned(26738, LDPC_TABLE_DATA_WIDTH)),
    246 => std_logic_vector(to_unsigned(6030, LDPC_TABLE_DATA_WIDTH)),
    247 => std_logic_vector(to_unsigned(505, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    248 => std_logic_vector(to_unsigned(85, LDPC_TABLE_DATA_WIDTH)),
    249 => std_logic_vector(to_unsigned(30326, LDPC_TABLE_DATA_WIDTH)),
    250 => std_logic_vector(to_unsigned(22298, LDPC_TABLE_DATA_WIDTH)),
    251 => std_logic_vector(to_unsigned(27562, LDPC_TABLE_DATA_WIDTH)),
    252 => std_logic_vector(to_unsigned(20131, LDPC_TABLE_DATA_WIDTH)),
    253 => std_logic_vector(to_unsigned(26390, LDPC_TABLE_DATA_WIDTH)),
    254 => std_logic_vector(to_unsigned(6247, LDPC_TABLE_DATA_WIDTH)),
    255 => std_logic_vector(to_unsigned(24791, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    256 => std_logic_vector(to_unsigned(86, LDPC_TABLE_DATA_WIDTH)),
    257 => std_logic_vector(to_unsigned(928, LDPC_TABLE_DATA_WIDTH)),
    258 => std_logic_vector(to_unsigned(29246, LDPC_TABLE_DATA_WIDTH)),
    259 => std_logic_vector(to_unsigned(21246, LDPC_TABLE_DATA_WIDTH)),
    260 => std_logic_vector(to_unsigned(12400, LDPC_TABLE_DATA_WIDTH)),
    261 => std_logic_vector(to_unsigned(15311, LDPC_TABLE_DATA_WIDTH)),
    262 => std_logic_vector(to_unsigned(32309, LDPC_TABLE_DATA_WIDTH)),
    263 => std_logic_vector(to_unsigned(18608, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    264 => std_logic_vector(to_unsigned(87, LDPC_TABLE_DATA_WIDTH)),
    265 => std_logic_vector(to_unsigned(20314, LDPC_TABLE_DATA_WIDTH)),
    266 => std_logic_vector(to_unsigned(6025, LDPC_TABLE_DATA_WIDTH)),
    267 => std_logic_vector(to_unsigned(26689, LDPC_TABLE_DATA_WIDTH)),
    268 => std_logic_vector(to_unsigned(16302, LDPC_TABLE_DATA_WIDTH)),
    269 => std_logic_vector(to_unsigned(2296, LDPC_TABLE_DATA_WIDTH)),
    270 => std_logic_vector(to_unsigned(3244, LDPC_TABLE_DATA_WIDTH)),
    271 => std_logic_vector(to_unsigned(19613, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    272 => std_logic_vector(to_unsigned(88, LDPC_TABLE_DATA_WIDTH)),
    273 => std_logic_vector(to_unsigned(6237, LDPC_TABLE_DATA_WIDTH)),
    274 => std_logic_vector(to_unsigned(11943, LDPC_TABLE_DATA_WIDTH)),
    275 => std_logic_vector(to_unsigned(22851, LDPC_TABLE_DATA_WIDTH)),
    276 => std_logic_vector(to_unsigned(15642, LDPC_TABLE_DATA_WIDTH)),
    277 => std_logic_vector(to_unsigned(23857, LDPC_TABLE_DATA_WIDTH)),
    278 => std_logic_vector(to_unsigned(15112, LDPC_TABLE_DATA_WIDTH)),
    279 => std_logic_vector(to_unsigned(20947, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    280 => std_logic_vector(to_unsigned(89, LDPC_TABLE_DATA_WIDTH)),
    281 => std_logic_vector(to_unsigned(26403, LDPC_TABLE_DATA_WIDTH)),
    282 => std_logic_vector(to_unsigned(25168, LDPC_TABLE_DATA_WIDTH)),
    283 => std_logic_vector(to_unsigned(19038, LDPC_TABLE_DATA_WIDTH)),
    284 => std_logic_vector(to_unsigned(18384, LDPC_TABLE_DATA_WIDTH)),
    285 => std_logic_vector(to_unsigned(8882, LDPC_TABLE_DATA_WIDTH)),
    286 => std_logic_vector(to_unsigned(12719, LDPC_TABLE_DATA_WIDTH)),
    287 => std_logic_vector(to_unsigned(7093, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    288 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    289 => std_logic_vector(to_unsigned(14567, LDPC_TABLE_DATA_WIDTH)),
    290 => std_logic_vector(to_unsigned(24965, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    291 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    292 => std_logic_vector(to_unsigned(3908, LDPC_TABLE_DATA_WIDTH)),
    293 => std_logic_vector(to_unsigned(100, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    294 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    295 => std_logic_vector(to_unsigned(10279, LDPC_TABLE_DATA_WIDTH)),
    296 => std_logic_vector(to_unsigned(240, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    297 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    298 => std_logic_vector(to_unsigned(24102, LDPC_TABLE_DATA_WIDTH)),
    299 => std_logic_vector(to_unsigned(764, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    300 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    301 => std_logic_vector(to_unsigned(12383, LDPC_TABLE_DATA_WIDTH)),
    302 => std_logic_vector(to_unsigned(4173, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    303 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    304 => std_logic_vector(to_unsigned(13861, LDPC_TABLE_DATA_WIDTH)),
    305 => std_logic_vector(to_unsigned(15918, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    306 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    307 => std_logic_vector(to_unsigned(21327, LDPC_TABLE_DATA_WIDTH)),
    308 => std_logic_vector(to_unsigned(1046, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    309 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    310 => std_logic_vector(to_unsigned(5288, LDPC_TABLE_DATA_WIDTH)),
    311 => std_logic_vector(to_unsigned(14579, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    312 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    313 => std_logic_vector(to_unsigned(28158, LDPC_TABLE_DATA_WIDTH)),
    314 => std_logic_vector(to_unsigned(8069, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    315 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    316 => std_logic_vector(to_unsigned(16583, LDPC_TABLE_DATA_WIDTH)),
    317 => std_logic_vector(to_unsigned(11098, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    318 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    319 => std_logic_vector(to_unsigned(16681, LDPC_TABLE_DATA_WIDTH)),
    320 => std_logic_vector(to_unsigned(28363, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    321 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    322 => std_logic_vector(to_unsigned(13980, LDPC_TABLE_DATA_WIDTH)),
    323 => std_logic_vector(to_unsigned(24725, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    324 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    325 => std_logic_vector(to_unsigned(32169, LDPC_TABLE_DATA_WIDTH)),
    326 => std_logic_vector(to_unsigned(17989, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    327 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    328 => std_logic_vector(to_unsigned(10907, LDPC_TABLE_DATA_WIDTH)),
    329 => std_logic_vector(to_unsigned(2767, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    330 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    331 => std_logic_vector(to_unsigned(21557, LDPC_TABLE_DATA_WIDTH)),
    332 => std_logic_vector(to_unsigned(3818, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    333 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    334 => std_logic_vector(to_unsigned(26676, LDPC_TABLE_DATA_WIDTH)),
    335 => std_logic_vector(to_unsigned(12422, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    336 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    337 => std_logic_vector(to_unsigned(7676, LDPC_TABLE_DATA_WIDTH)),
    338 => std_logic_vector(to_unsigned(8754, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    339 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    340 => std_logic_vector(to_unsigned(14905, LDPC_TABLE_DATA_WIDTH)),
    341 => std_logic_vector(to_unsigned(20232, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    342 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    343 => std_logic_vector(to_unsigned(15719, LDPC_TABLE_DATA_WIDTH)),
    344 => std_logic_vector(to_unsigned(24646, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    345 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    346 => std_logic_vector(to_unsigned(31942, LDPC_TABLE_DATA_WIDTH)),
    347 => std_logic_vector(to_unsigned(8589, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    348 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    349 => std_logic_vector(to_unsigned(19978, LDPC_TABLE_DATA_WIDTH)),
    350 => std_logic_vector(to_unsigned(27197, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    351 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    352 => std_logic_vector(to_unsigned(27060, LDPC_TABLE_DATA_WIDTH)),
    353 => std_logic_vector(to_unsigned(15071, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    354 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    355 => std_logic_vector(to_unsigned(6071, LDPC_TABLE_DATA_WIDTH)),
    356 => std_logic_vector(to_unsigned(26649, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    357 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    358 => std_logic_vector(to_unsigned(10393, LDPC_TABLE_DATA_WIDTH)),
    359 => std_logic_vector(to_unsigned(11176, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    360 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    361 => std_logic_vector(to_unsigned(9597, LDPC_TABLE_DATA_WIDTH)),
    362 => std_logic_vector(to_unsigned(13370, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    363 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    364 => std_logic_vector(to_unsigned(7081, LDPC_TABLE_DATA_WIDTH)),
    365 => std_logic_vector(to_unsigned(17677, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    366 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    367 => std_logic_vector(to_unsigned(1433, LDPC_TABLE_DATA_WIDTH)),
    368 => std_logic_vector(to_unsigned(19513, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    369 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    370 => std_logic_vector(to_unsigned(26925, LDPC_TABLE_DATA_WIDTH)),
    371 => std_logic_vector(to_unsigned(9014, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    372 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    373 => std_logic_vector(to_unsigned(19202, LDPC_TABLE_DATA_WIDTH)),
    374 => std_logic_vector(to_unsigned(8900, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    375 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    376 => std_logic_vector(to_unsigned(18152, LDPC_TABLE_DATA_WIDTH)),
    377 => std_logic_vector(to_unsigned(30647, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    378 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    379 => std_logic_vector(to_unsigned(20803, LDPC_TABLE_DATA_WIDTH)),
    380 => std_logic_vector(to_unsigned(1737, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    381 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    382 => std_logic_vector(to_unsigned(11804, LDPC_TABLE_DATA_WIDTH)),
    383 => std_logic_vector(to_unsigned(25221, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    384 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    385 => std_logic_vector(to_unsigned(31683, LDPC_TABLE_DATA_WIDTH)),
    386 => std_logic_vector(to_unsigned(17783, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    387 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    388 => std_logic_vector(to_unsigned(29694, LDPC_TABLE_DATA_WIDTH)),
    389 => std_logic_vector(to_unsigned(9345, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    390 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    391 => std_logic_vector(to_unsigned(12280, LDPC_TABLE_DATA_WIDTH)),
    392 => std_logic_vector(to_unsigned(26611, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    393 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    394 => std_logic_vector(to_unsigned(6526, LDPC_TABLE_DATA_WIDTH)),
    395 => std_logic_vector(to_unsigned(26122, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    396 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    397 => std_logic_vector(to_unsigned(26165, LDPC_TABLE_DATA_WIDTH)),
    398 => std_logic_vector(to_unsigned(11241, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    399 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    400 => std_logic_vector(to_unsigned(7666, LDPC_TABLE_DATA_WIDTH)),
    401 => std_logic_vector(to_unsigned(26962, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    402 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    403 => std_logic_vector(to_unsigned(16290, LDPC_TABLE_DATA_WIDTH)),
    404 => std_logic_vector(to_unsigned(8480, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    405 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    406 => std_logic_vector(to_unsigned(11774, LDPC_TABLE_DATA_WIDTH)),
    407 => std_logic_vector(to_unsigned(10120, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    408 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    409 => std_logic_vector(to_unsigned(30051, LDPC_TABLE_DATA_WIDTH)),
    410 => std_logic_vector(to_unsigned(30426, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    411 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    412 => std_logic_vector(to_unsigned(1335, LDPC_TABLE_DATA_WIDTH)),
    413 => std_logic_vector(to_unsigned(15424, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    414 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    415 => std_logic_vector(to_unsigned(6865, LDPC_TABLE_DATA_WIDTH)),
    416 => std_logic_vector(to_unsigned(17742, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    417 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    418 => std_logic_vector(to_unsigned(31779, LDPC_TABLE_DATA_WIDTH)),
    419 => std_logic_vector(to_unsigned(12489, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    420 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    421 => std_logic_vector(to_unsigned(32120, LDPC_TABLE_DATA_WIDTH)),
    422 => std_logic_vector(to_unsigned(21001, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    423 => std_logic_vector(to_unsigned(45, LDPC_TABLE_DATA_WIDTH)),
    424 => std_logic_vector(to_unsigned(14508, LDPC_TABLE_DATA_WIDTH)),
    425 => std_logic_vector(to_unsigned(6996, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    426 => std_logic_vector(to_unsigned(46, LDPC_TABLE_DATA_WIDTH)),
    427 => std_logic_vector(to_unsigned(979, LDPC_TABLE_DATA_WIDTH)),
    428 => std_logic_vector(to_unsigned(25024, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    429 => std_logic_vector(to_unsigned(47, LDPC_TABLE_DATA_WIDTH)),
    430 => std_logic_vector(to_unsigned(4554, LDPC_TABLE_DATA_WIDTH)),
    431 => std_logic_vector(to_unsigned(21896, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    432 => std_logic_vector(to_unsigned(48, LDPC_TABLE_DATA_WIDTH)),
    433 => std_logic_vector(to_unsigned(7989, LDPC_TABLE_DATA_WIDTH)),
    434 => std_logic_vector(to_unsigned(21777, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    435 => std_logic_vector(to_unsigned(49, LDPC_TABLE_DATA_WIDTH)),
    436 => std_logic_vector(to_unsigned(4972, LDPC_TABLE_DATA_WIDTH)),
    437 => std_logic_vector(to_unsigned(20661, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    438 => std_logic_vector(to_unsigned(50, LDPC_TABLE_DATA_WIDTH)),
    439 => std_logic_vector(to_unsigned(6612, LDPC_TABLE_DATA_WIDTH)),
    440 => std_logic_vector(to_unsigned(2730, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    441 => std_logic_vector(to_unsigned(51, LDPC_TABLE_DATA_WIDTH)),
    442 => std_logic_vector(to_unsigned(12742, LDPC_TABLE_DATA_WIDTH)),
    443 => std_logic_vector(to_unsigned(4418, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    444 => std_logic_vector(to_unsigned(52, LDPC_TABLE_DATA_WIDTH)),
    445 => std_logic_vector(to_unsigned(29194, LDPC_TABLE_DATA_WIDTH)),
    446 => std_logic_vector(to_unsigned(595, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    447 => std_logic_vector(to_unsigned(53, LDPC_TABLE_DATA_WIDTH)),
    448 => std_logic_vector(to_unsigned(19267, LDPC_TABLE_DATA_WIDTH)),
    449 => std_logic_vector(to_unsigned(20113, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C1_3
    450 => std_logic_vector(to_unsigned(34903, LDPC_TABLE_DATA_WIDTH)),
    451 => std_logic_vector(to_unsigned(20927, LDPC_TABLE_DATA_WIDTH)),
    452 => std_logic_vector(to_unsigned(32093, LDPC_TABLE_DATA_WIDTH)),
    453 => std_logic_vector(to_unsigned(1052, LDPC_TABLE_DATA_WIDTH)),
    454 => std_logic_vector(to_unsigned(25611, LDPC_TABLE_DATA_WIDTH)),
    455 => std_logic_vector(to_unsigned(16093, LDPC_TABLE_DATA_WIDTH)),
    456 => std_logic_vector(to_unsigned(16454, LDPC_TABLE_DATA_WIDTH)),
    457 => std_logic_vector(to_unsigned(5520, LDPC_TABLE_DATA_WIDTH)),
    458 => std_logic_vector(to_unsigned(506, LDPC_TABLE_DATA_WIDTH)),
    459 => std_logic_vector(to_unsigned(37399, LDPC_TABLE_DATA_WIDTH)),
    460 => std_logic_vector(to_unsigned(18518, LDPC_TABLE_DATA_WIDTH)),
    461 => std_logic_vector(to_unsigned(21120, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    462 => std_logic_vector(to_unsigned(11636, LDPC_TABLE_DATA_WIDTH)),
    463 => std_logic_vector(to_unsigned(14594, LDPC_TABLE_DATA_WIDTH)),
    464 => std_logic_vector(to_unsigned(22158, LDPC_TABLE_DATA_WIDTH)),
    465 => std_logic_vector(to_unsigned(14763, LDPC_TABLE_DATA_WIDTH)),
    466 => std_logic_vector(to_unsigned(15333, LDPC_TABLE_DATA_WIDTH)),
    467 => std_logic_vector(to_unsigned(6838, LDPC_TABLE_DATA_WIDTH)),
    468 => std_logic_vector(to_unsigned(22222, LDPC_TABLE_DATA_WIDTH)),
    469 => std_logic_vector(to_unsigned(37856, LDPC_TABLE_DATA_WIDTH)),
    470 => std_logic_vector(to_unsigned(14985, LDPC_TABLE_DATA_WIDTH)),
    471 => std_logic_vector(to_unsigned(31041, LDPC_TABLE_DATA_WIDTH)),
    472 => std_logic_vector(to_unsigned(18704, LDPC_TABLE_DATA_WIDTH)),
    473 => std_logic_vector(to_unsigned(32910, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    474 => std_logic_vector(to_unsigned(17449, LDPC_TABLE_DATA_WIDTH)),
    475 => std_logic_vector(to_unsigned(1665, LDPC_TABLE_DATA_WIDTH)),
    476 => std_logic_vector(to_unsigned(35639, LDPC_TABLE_DATA_WIDTH)),
    477 => std_logic_vector(to_unsigned(16624, LDPC_TABLE_DATA_WIDTH)),
    478 => std_logic_vector(to_unsigned(12867, LDPC_TABLE_DATA_WIDTH)),
    479 => std_logic_vector(to_unsigned(12449, LDPC_TABLE_DATA_WIDTH)),
    480 => std_logic_vector(to_unsigned(10241, LDPC_TABLE_DATA_WIDTH)),
    481 => std_logic_vector(to_unsigned(11650, LDPC_TABLE_DATA_WIDTH)),
    482 => std_logic_vector(to_unsigned(25622, LDPC_TABLE_DATA_WIDTH)),
    483 => std_logic_vector(to_unsigned(34372, LDPC_TABLE_DATA_WIDTH)),
    484 => std_logic_vector(to_unsigned(19878, LDPC_TABLE_DATA_WIDTH)),
    485 => std_logic_vector(to_unsigned(26894, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    486 => std_logic_vector(to_unsigned(29235, LDPC_TABLE_DATA_WIDTH)),
    487 => std_logic_vector(to_unsigned(19780, LDPC_TABLE_DATA_WIDTH)),
    488 => std_logic_vector(to_unsigned(36056, LDPC_TABLE_DATA_WIDTH)),
    489 => std_logic_vector(to_unsigned(20129, LDPC_TABLE_DATA_WIDTH)),
    490 => std_logic_vector(to_unsigned(20029, LDPC_TABLE_DATA_WIDTH)),
    491 => std_logic_vector(to_unsigned(5457, LDPC_TABLE_DATA_WIDTH)),
    492 => std_logic_vector(to_unsigned(8157, LDPC_TABLE_DATA_WIDTH)),
    493 => std_logic_vector(to_unsigned(35554, LDPC_TABLE_DATA_WIDTH)),
    494 => std_logic_vector(to_unsigned(21237, LDPC_TABLE_DATA_WIDTH)),
    495 => std_logic_vector(to_unsigned(7943, LDPC_TABLE_DATA_WIDTH)),
    496 => std_logic_vector(to_unsigned(13873, LDPC_TABLE_DATA_WIDTH)),
    497 => std_logic_vector(to_unsigned(14980, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    498 => std_logic_vector(to_unsigned(9912, LDPC_TABLE_DATA_WIDTH)),
    499 => std_logic_vector(to_unsigned(7143, LDPC_TABLE_DATA_WIDTH)),
    500 => std_logic_vector(to_unsigned(35911, LDPC_TABLE_DATA_WIDTH)),
    501 => std_logic_vector(to_unsigned(12043, LDPC_TABLE_DATA_WIDTH)),
    502 => std_logic_vector(to_unsigned(17360, LDPC_TABLE_DATA_WIDTH)),
    503 => std_logic_vector(to_unsigned(37253, LDPC_TABLE_DATA_WIDTH)),
    504 => std_logic_vector(to_unsigned(25588, LDPC_TABLE_DATA_WIDTH)),
    505 => std_logic_vector(to_unsigned(11827, LDPC_TABLE_DATA_WIDTH)),
    506 => std_logic_vector(to_unsigned(29152, LDPC_TABLE_DATA_WIDTH)),
    507 => std_logic_vector(to_unsigned(21936, LDPC_TABLE_DATA_WIDTH)),
    508 => std_logic_vector(to_unsigned(24125, LDPC_TABLE_DATA_WIDTH)),
    509 => std_logic_vector(to_unsigned(40870, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    510 => std_logic_vector(to_unsigned(40701, LDPC_TABLE_DATA_WIDTH)),
    511 => std_logic_vector(to_unsigned(36035, LDPC_TABLE_DATA_WIDTH)),
    512 => std_logic_vector(to_unsigned(39556, LDPC_TABLE_DATA_WIDTH)),
    513 => std_logic_vector(to_unsigned(12366, LDPC_TABLE_DATA_WIDTH)),
    514 => std_logic_vector(to_unsigned(19946, LDPC_TABLE_DATA_WIDTH)),
    515 => std_logic_vector(to_unsigned(29072, LDPC_TABLE_DATA_WIDTH)),
    516 => std_logic_vector(to_unsigned(16365, LDPC_TABLE_DATA_WIDTH)),
    517 => std_logic_vector(to_unsigned(35495, LDPC_TABLE_DATA_WIDTH)),
    518 => std_logic_vector(to_unsigned(22686, LDPC_TABLE_DATA_WIDTH)),
    519 => std_logic_vector(to_unsigned(11106, LDPC_TABLE_DATA_WIDTH)),
    520 => std_logic_vector(to_unsigned(8756, LDPC_TABLE_DATA_WIDTH)),
    521 => std_logic_vector(to_unsigned(34863, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    522 => std_logic_vector(to_unsigned(19165, LDPC_TABLE_DATA_WIDTH)),
    523 => std_logic_vector(to_unsigned(15702, LDPC_TABLE_DATA_WIDTH)),
    524 => std_logic_vector(to_unsigned(13536, LDPC_TABLE_DATA_WIDTH)),
    525 => std_logic_vector(to_unsigned(40238, LDPC_TABLE_DATA_WIDTH)),
    526 => std_logic_vector(to_unsigned(4465, LDPC_TABLE_DATA_WIDTH)),
    527 => std_logic_vector(to_unsigned(40034, LDPC_TABLE_DATA_WIDTH)),
    528 => std_logic_vector(to_unsigned(40590, LDPC_TABLE_DATA_WIDTH)),
    529 => std_logic_vector(to_unsigned(37540, LDPC_TABLE_DATA_WIDTH)),
    530 => std_logic_vector(to_unsigned(17162, LDPC_TABLE_DATA_WIDTH)),
    531 => std_logic_vector(to_unsigned(1712, LDPC_TABLE_DATA_WIDTH)),
    532 => std_logic_vector(to_unsigned(20577, LDPC_TABLE_DATA_WIDTH)),
    533 => std_logic_vector(to_unsigned(14138, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    534 => std_logic_vector(to_unsigned(31338, LDPC_TABLE_DATA_WIDTH)),
    535 => std_logic_vector(to_unsigned(19342, LDPC_TABLE_DATA_WIDTH)),
    536 => std_logic_vector(to_unsigned(9301, LDPC_TABLE_DATA_WIDTH)),
    537 => std_logic_vector(to_unsigned(39375, LDPC_TABLE_DATA_WIDTH)),
    538 => std_logic_vector(to_unsigned(3211, LDPC_TABLE_DATA_WIDTH)),
    539 => std_logic_vector(to_unsigned(1316, LDPC_TABLE_DATA_WIDTH)),
    540 => std_logic_vector(to_unsigned(33409, LDPC_TABLE_DATA_WIDTH)),
    541 => std_logic_vector(to_unsigned(28670, LDPC_TABLE_DATA_WIDTH)),
    542 => std_logic_vector(to_unsigned(12282, LDPC_TABLE_DATA_WIDTH)),
    543 => std_logic_vector(to_unsigned(6118, LDPC_TABLE_DATA_WIDTH)),
    544 => std_logic_vector(to_unsigned(29236, LDPC_TABLE_DATA_WIDTH)),
    545 => std_logic_vector(to_unsigned(35787, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    546 => std_logic_vector(to_unsigned(11504, LDPC_TABLE_DATA_WIDTH)),
    547 => std_logic_vector(to_unsigned(30506, LDPC_TABLE_DATA_WIDTH)),
    548 => std_logic_vector(to_unsigned(19558, LDPC_TABLE_DATA_WIDTH)),
    549 => std_logic_vector(to_unsigned(5100, LDPC_TABLE_DATA_WIDTH)),
    550 => std_logic_vector(to_unsigned(24188, LDPC_TABLE_DATA_WIDTH)),
    551 => std_logic_vector(to_unsigned(24738, LDPC_TABLE_DATA_WIDTH)),
    552 => std_logic_vector(to_unsigned(30397, LDPC_TABLE_DATA_WIDTH)),
    553 => std_logic_vector(to_unsigned(33775, LDPC_TABLE_DATA_WIDTH)),
    554 => std_logic_vector(to_unsigned(9699, LDPC_TABLE_DATA_WIDTH)),
    555 => std_logic_vector(to_unsigned(6215, LDPC_TABLE_DATA_WIDTH)),
    556 => std_logic_vector(to_unsigned(3397, LDPC_TABLE_DATA_WIDTH)),
    557 => std_logic_vector(to_unsigned(37451, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    558 => std_logic_vector(to_unsigned(34689, LDPC_TABLE_DATA_WIDTH)),
    559 => std_logic_vector(to_unsigned(23126, LDPC_TABLE_DATA_WIDTH)),
    560 => std_logic_vector(to_unsigned(7571, LDPC_TABLE_DATA_WIDTH)),
    561 => std_logic_vector(to_unsigned(1058, LDPC_TABLE_DATA_WIDTH)),
    562 => std_logic_vector(to_unsigned(12127, LDPC_TABLE_DATA_WIDTH)),
    563 => std_logic_vector(to_unsigned(27518, LDPC_TABLE_DATA_WIDTH)),
    564 => std_logic_vector(to_unsigned(23064, LDPC_TABLE_DATA_WIDTH)),
    565 => std_logic_vector(to_unsigned(11265, LDPC_TABLE_DATA_WIDTH)),
    566 => std_logic_vector(to_unsigned(14867, LDPC_TABLE_DATA_WIDTH)),
    567 => std_logic_vector(to_unsigned(30451, LDPC_TABLE_DATA_WIDTH)),
    568 => std_logic_vector(to_unsigned(28289, LDPC_TABLE_DATA_WIDTH)),
    569 => std_logic_vector(to_unsigned(2966, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    570 => std_logic_vector(to_unsigned(11660, LDPC_TABLE_DATA_WIDTH)),
    571 => std_logic_vector(to_unsigned(15334, LDPC_TABLE_DATA_WIDTH)),
    572 => std_logic_vector(to_unsigned(16867, LDPC_TABLE_DATA_WIDTH)),
    573 => std_logic_vector(to_unsigned(15160, LDPC_TABLE_DATA_WIDTH)),
    574 => std_logic_vector(to_unsigned(38343, LDPC_TABLE_DATA_WIDTH)),
    575 => std_logic_vector(to_unsigned(3778, LDPC_TABLE_DATA_WIDTH)),
    576 => std_logic_vector(to_unsigned(4265, LDPC_TABLE_DATA_WIDTH)),
    577 => std_logic_vector(to_unsigned(39139, LDPC_TABLE_DATA_WIDTH)),
    578 => std_logic_vector(to_unsigned(17293, LDPC_TABLE_DATA_WIDTH)),
    579 => std_logic_vector(to_unsigned(26229, LDPC_TABLE_DATA_WIDTH)),
    580 => std_logic_vector(to_unsigned(42604, LDPC_TABLE_DATA_WIDTH)),
    581 => std_logic_vector(to_unsigned(13486, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    582 => std_logic_vector(to_unsigned(31497, LDPC_TABLE_DATA_WIDTH)),
    583 => std_logic_vector(to_unsigned(1365, LDPC_TABLE_DATA_WIDTH)),
    584 => std_logic_vector(to_unsigned(14828, LDPC_TABLE_DATA_WIDTH)),
    585 => std_logic_vector(to_unsigned(7453, LDPC_TABLE_DATA_WIDTH)),
    586 => std_logic_vector(to_unsigned(26350, LDPC_TABLE_DATA_WIDTH)),
    587 => std_logic_vector(to_unsigned(41346, LDPC_TABLE_DATA_WIDTH)),
    588 => std_logic_vector(to_unsigned(28643, LDPC_TABLE_DATA_WIDTH)),
    589 => std_logic_vector(to_unsigned(23421, LDPC_TABLE_DATA_WIDTH)),
    590 => std_logic_vector(to_unsigned(8354, LDPC_TABLE_DATA_WIDTH)),
    591 => std_logic_vector(to_unsigned(16255, LDPC_TABLE_DATA_WIDTH)),
    592 => std_logic_vector(to_unsigned(11055, LDPC_TABLE_DATA_WIDTH)),
    593 => std_logic_vector(to_unsigned(24279, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    594 => std_logic_vector(to_unsigned(15687, LDPC_TABLE_DATA_WIDTH)),
    595 => std_logic_vector(to_unsigned(12467, LDPC_TABLE_DATA_WIDTH)),
    596 => std_logic_vector(to_unsigned(13906, LDPC_TABLE_DATA_WIDTH)),
    597 => std_logic_vector(to_unsigned(5215, LDPC_TABLE_DATA_WIDTH)),
    598 => std_logic_vector(to_unsigned(41328, LDPC_TABLE_DATA_WIDTH)),
    599 => std_logic_vector(to_unsigned(23755, LDPC_TABLE_DATA_WIDTH)),
    600 => std_logic_vector(to_unsigned(20800, LDPC_TABLE_DATA_WIDTH)),
    601 => std_logic_vector(to_unsigned(6447, LDPC_TABLE_DATA_WIDTH)),
    602 => std_logic_vector(to_unsigned(7970, LDPC_TABLE_DATA_WIDTH)),
    603 => std_logic_vector(to_unsigned(2803, LDPC_TABLE_DATA_WIDTH)),
    604 => std_logic_vector(to_unsigned(33262, LDPC_TABLE_DATA_WIDTH)),
    605 => std_logic_vector(to_unsigned(39843, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    606 => std_logic_vector(to_unsigned(5363, LDPC_TABLE_DATA_WIDTH)),
    607 => std_logic_vector(to_unsigned(22469, LDPC_TABLE_DATA_WIDTH)),
    608 => std_logic_vector(to_unsigned(38091, LDPC_TABLE_DATA_WIDTH)),
    609 => std_logic_vector(to_unsigned(28457, LDPC_TABLE_DATA_WIDTH)),
    610 => std_logic_vector(to_unsigned(36696, LDPC_TABLE_DATA_WIDTH)),
    611 => std_logic_vector(to_unsigned(34471, LDPC_TABLE_DATA_WIDTH)),
    612 => std_logic_vector(to_unsigned(23619, LDPC_TABLE_DATA_WIDTH)),
    613 => std_logic_vector(to_unsigned(2404, LDPC_TABLE_DATA_WIDTH)),
    614 => std_logic_vector(to_unsigned(24229, LDPC_TABLE_DATA_WIDTH)),
    615 => std_logic_vector(to_unsigned(41754, LDPC_TABLE_DATA_WIDTH)),
    616 => std_logic_vector(to_unsigned(1297, LDPC_TABLE_DATA_WIDTH)),
    617 => std_logic_vector(to_unsigned(18563, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    618 => std_logic_vector(to_unsigned(3673, LDPC_TABLE_DATA_WIDTH)),
    619 => std_logic_vector(to_unsigned(39070, LDPC_TABLE_DATA_WIDTH)),
    620 => std_logic_vector(to_unsigned(14480, LDPC_TABLE_DATA_WIDTH)),
    621 => std_logic_vector(to_unsigned(30279, LDPC_TABLE_DATA_WIDTH)),
    622 => std_logic_vector(to_unsigned(37483, LDPC_TABLE_DATA_WIDTH)),
    623 => std_logic_vector(to_unsigned(7580, LDPC_TABLE_DATA_WIDTH)),
    624 => std_logic_vector(to_unsigned(29519, LDPC_TABLE_DATA_WIDTH)),
    625 => std_logic_vector(to_unsigned(30519, LDPC_TABLE_DATA_WIDTH)),
    626 => std_logic_vector(to_unsigned(39831, LDPC_TABLE_DATA_WIDTH)),
    627 => std_logic_vector(to_unsigned(20252, LDPC_TABLE_DATA_WIDTH)),
    628 => std_logic_vector(to_unsigned(18132, LDPC_TABLE_DATA_WIDTH)),
    629 => std_logic_vector(to_unsigned(20010, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    630 => std_logic_vector(to_unsigned(34386, LDPC_TABLE_DATA_WIDTH)),
    631 => std_logic_vector(to_unsigned(7252, LDPC_TABLE_DATA_WIDTH)),
    632 => std_logic_vector(to_unsigned(27526, LDPC_TABLE_DATA_WIDTH)),
    633 => std_logic_vector(to_unsigned(12950, LDPC_TABLE_DATA_WIDTH)),
    634 => std_logic_vector(to_unsigned(6875, LDPC_TABLE_DATA_WIDTH)),
    635 => std_logic_vector(to_unsigned(43020, LDPC_TABLE_DATA_WIDTH)),
    636 => std_logic_vector(to_unsigned(31566, LDPC_TABLE_DATA_WIDTH)),
    637 => std_logic_vector(to_unsigned(39069, LDPC_TABLE_DATA_WIDTH)),
    638 => std_logic_vector(to_unsigned(18985, LDPC_TABLE_DATA_WIDTH)),
    639 => std_logic_vector(to_unsigned(15541, LDPC_TABLE_DATA_WIDTH)),
    640 => std_logic_vector(to_unsigned(40020, LDPC_TABLE_DATA_WIDTH)),
    641 => std_logic_vector(to_unsigned(16715, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    642 => std_logic_vector(to_unsigned(1721, LDPC_TABLE_DATA_WIDTH)),
    643 => std_logic_vector(to_unsigned(37332, LDPC_TABLE_DATA_WIDTH)),
    644 => std_logic_vector(to_unsigned(39953, LDPC_TABLE_DATA_WIDTH)),
    645 => std_logic_vector(to_unsigned(17430, LDPC_TABLE_DATA_WIDTH)),
    646 => std_logic_vector(to_unsigned(32134, LDPC_TABLE_DATA_WIDTH)),
    647 => std_logic_vector(to_unsigned(29162, LDPC_TABLE_DATA_WIDTH)),
    648 => std_logic_vector(to_unsigned(10490, LDPC_TABLE_DATA_WIDTH)),
    649 => std_logic_vector(to_unsigned(12971, LDPC_TABLE_DATA_WIDTH)),
    650 => std_logic_vector(to_unsigned(28581, LDPC_TABLE_DATA_WIDTH)),
    651 => std_logic_vector(to_unsigned(29331, LDPC_TABLE_DATA_WIDTH)),
    652 => std_logic_vector(to_unsigned(6489, LDPC_TABLE_DATA_WIDTH)),
    653 => std_logic_vector(to_unsigned(35383, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    654 => std_logic_vector(to_unsigned(736, LDPC_TABLE_DATA_WIDTH)),
    655 => std_logic_vector(to_unsigned(7022, LDPC_TABLE_DATA_WIDTH)),
    656 => std_logic_vector(to_unsigned(42349, LDPC_TABLE_DATA_WIDTH)),
    657 => std_logic_vector(to_unsigned(8783, LDPC_TABLE_DATA_WIDTH)),
    658 => std_logic_vector(to_unsigned(6767, LDPC_TABLE_DATA_WIDTH)),
    659 => std_logic_vector(to_unsigned(11871, LDPC_TABLE_DATA_WIDTH)),
    660 => std_logic_vector(to_unsigned(21675, LDPC_TABLE_DATA_WIDTH)),
    661 => std_logic_vector(to_unsigned(10325, LDPC_TABLE_DATA_WIDTH)),
    662 => std_logic_vector(to_unsigned(11548, LDPC_TABLE_DATA_WIDTH)),
    663 => std_logic_vector(to_unsigned(25978, LDPC_TABLE_DATA_WIDTH)),
    664 => std_logic_vector(to_unsigned(431, LDPC_TABLE_DATA_WIDTH)),
    665 => std_logic_vector(to_unsigned(24085, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    666 => std_logic_vector(to_unsigned(1925, LDPC_TABLE_DATA_WIDTH)),
    667 => std_logic_vector(to_unsigned(10602, LDPC_TABLE_DATA_WIDTH)),
    668 => std_logic_vector(to_unsigned(28585, LDPC_TABLE_DATA_WIDTH)),
    669 => std_logic_vector(to_unsigned(12170, LDPC_TABLE_DATA_WIDTH)),
    670 => std_logic_vector(to_unsigned(15156, LDPC_TABLE_DATA_WIDTH)),
    671 => std_logic_vector(to_unsigned(34404, LDPC_TABLE_DATA_WIDTH)),
    672 => std_logic_vector(to_unsigned(8351, LDPC_TABLE_DATA_WIDTH)),
    673 => std_logic_vector(to_unsigned(13273, LDPC_TABLE_DATA_WIDTH)),
    674 => std_logic_vector(to_unsigned(20208, LDPC_TABLE_DATA_WIDTH)),
    675 => std_logic_vector(to_unsigned(5800, LDPC_TABLE_DATA_WIDTH)),
    676 => std_logic_vector(to_unsigned(15367, LDPC_TABLE_DATA_WIDTH)),
    677 => std_logic_vector(to_unsigned(21764, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    678 => std_logic_vector(to_unsigned(16279, LDPC_TABLE_DATA_WIDTH)),
    679 => std_logic_vector(to_unsigned(37832, LDPC_TABLE_DATA_WIDTH)),
    680 => std_logic_vector(to_unsigned(34792, LDPC_TABLE_DATA_WIDTH)),
    681 => std_logic_vector(to_unsigned(21250, LDPC_TABLE_DATA_WIDTH)),
    682 => std_logic_vector(to_unsigned(34192, LDPC_TABLE_DATA_WIDTH)),
    683 => std_logic_vector(to_unsigned(7406, LDPC_TABLE_DATA_WIDTH)),
    684 => std_logic_vector(to_unsigned(41488, LDPC_TABLE_DATA_WIDTH)),
    685 => std_logic_vector(to_unsigned(18346, LDPC_TABLE_DATA_WIDTH)),
    686 => std_logic_vector(to_unsigned(29227, LDPC_TABLE_DATA_WIDTH)),
    687 => std_logic_vector(to_unsigned(26127, LDPC_TABLE_DATA_WIDTH)),
    688 => std_logic_vector(to_unsigned(25493, LDPC_TABLE_DATA_WIDTH)),
    689 => std_logic_vector(to_unsigned(7048, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    690 => std_logic_vector(to_unsigned(39948, LDPC_TABLE_DATA_WIDTH)),
    691 => std_logic_vector(to_unsigned(28229, LDPC_TABLE_DATA_WIDTH)),
    692 => std_logic_vector(to_unsigned(24899, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    693 => std_logic_vector(to_unsigned(17408, LDPC_TABLE_DATA_WIDTH)),
    694 => std_logic_vector(to_unsigned(14274, LDPC_TABLE_DATA_WIDTH)),
    695 => std_logic_vector(to_unsigned(38993, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    696 => std_logic_vector(to_unsigned(38774, LDPC_TABLE_DATA_WIDTH)),
    697 => std_logic_vector(to_unsigned(15968, LDPC_TABLE_DATA_WIDTH)),
    698 => std_logic_vector(to_unsigned(28459, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    699 => std_logic_vector(to_unsigned(41404, LDPC_TABLE_DATA_WIDTH)),
    700 => std_logic_vector(to_unsigned(27249, LDPC_TABLE_DATA_WIDTH)),
    701 => std_logic_vector(to_unsigned(27425, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    702 => std_logic_vector(to_unsigned(41229, LDPC_TABLE_DATA_WIDTH)),
    703 => std_logic_vector(to_unsigned(6082, LDPC_TABLE_DATA_WIDTH)),
    704 => std_logic_vector(to_unsigned(43114, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    705 => std_logic_vector(to_unsigned(13957, LDPC_TABLE_DATA_WIDTH)),
    706 => std_logic_vector(to_unsigned(4979, LDPC_TABLE_DATA_WIDTH)),
    707 => std_logic_vector(to_unsigned(40654, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    708 => std_logic_vector(to_unsigned(3093, LDPC_TABLE_DATA_WIDTH)),
    709 => std_logic_vector(to_unsigned(3438, LDPC_TABLE_DATA_WIDTH)),
    710 => std_logic_vector(to_unsigned(34992, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    711 => std_logic_vector(to_unsigned(34082, LDPC_TABLE_DATA_WIDTH)),
    712 => std_logic_vector(to_unsigned(6172, LDPC_TABLE_DATA_WIDTH)),
    713 => std_logic_vector(to_unsigned(28760, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    714 => std_logic_vector(to_unsigned(42210, LDPC_TABLE_DATA_WIDTH)),
    715 => std_logic_vector(to_unsigned(34141, LDPC_TABLE_DATA_WIDTH)),
    716 => std_logic_vector(to_unsigned(41021, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    717 => std_logic_vector(to_unsigned(14705, LDPC_TABLE_DATA_WIDTH)),
    718 => std_logic_vector(to_unsigned(17783, LDPC_TABLE_DATA_WIDTH)),
    719 => std_logic_vector(to_unsigned(10134, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    720 => std_logic_vector(to_unsigned(41755, LDPC_TABLE_DATA_WIDTH)),
    721 => std_logic_vector(to_unsigned(39884, LDPC_TABLE_DATA_WIDTH)),
    722 => std_logic_vector(to_unsigned(22773, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    723 => std_logic_vector(to_unsigned(14615, LDPC_TABLE_DATA_WIDTH)),
    724 => std_logic_vector(to_unsigned(15593, LDPC_TABLE_DATA_WIDTH)),
    725 => std_logic_vector(to_unsigned(1642, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    726 => std_logic_vector(to_unsigned(29111, LDPC_TABLE_DATA_WIDTH)),
    727 => std_logic_vector(to_unsigned(37061, LDPC_TABLE_DATA_WIDTH)),
    728 => std_logic_vector(to_unsigned(39860, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    729 => std_logic_vector(to_unsigned(9579, LDPC_TABLE_DATA_WIDTH)),
    730 => std_logic_vector(to_unsigned(33552, LDPC_TABLE_DATA_WIDTH)),
    731 => std_logic_vector(to_unsigned(633, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    732 => std_logic_vector(to_unsigned(12951, LDPC_TABLE_DATA_WIDTH)),
    733 => std_logic_vector(to_unsigned(21137, LDPC_TABLE_DATA_WIDTH)),
    734 => std_logic_vector(to_unsigned(39608, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    735 => std_logic_vector(to_unsigned(38244, LDPC_TABLE_DATA_WIDTH)),
    736 => std_logic_vector(to_unsigned(27361, LDPC_TABLE_DATA_WIDTH)),
    737 => std_logic_vector(to_unsigned(29417, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    738 => std_logic_vector(to_unsigned(2939, LDPC_TABLE_DATA_WIDTH)),
    739 => std_logic_vector(to_unsigned(10172, LDPC_TABLE_DATA_WIDTH)),
    740 => std_logic_vector(to_unsigned(36479, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    741 => std_logic_vector(to_unsigned(29094, LDPC_TABLE_DATA_WIDTH)),
    742 => std_logic_vector(to_unsigned(5357, LDPC_TABLE_DATA_WIDTH)),
    743 => std_logic_vector(to_unsigned(19224, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    744 => std_logic_vector(to_unsigned(9562, LDPC_TABLE_DATA_WIDTH)),
    745 => std_logic_vector(to_unsigned(24436, LDPC_TABLE_DATA_WIDTH)),
    746 => std_logic_vector(to_unsigned(28637, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    747 => std_logic_vector(to_unsigned(40177, LDPC_TABLE_DATA_WIDTH)),
    748 => std_logic_vector(to_unsigned(2326, LDPC_TABLE_DATA_WIDTH)),
    749 => std_logic_vector(to_unsigned(13504, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    750 => std_logic_vector(to_unsigned(6834, LDPC_TABLE_DATA_WIDTH)),
    751 => std_logic_vector(to_unsigned(21583, LDPC_TABLE_DATA_WIDTH)),
    752 => std_logic_vector(to_unsigned(42516, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    753 => std_logic_vector(to_unsigned(40651, LDPC_TABLE_DATA_WIDTH)),
    754 => std_logic_vector(to_unsigned(42810, LDPC_TABLE_DATA_WIDTH)),
    755 => std_logic_vector(to_unsigned(25709, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    756 => std_logic_vector(to_unsigned(31557, LDPC_TABLE_DATA_WIDTH)),
    757 => std_logic_vector(to_unsigned(32138, LDPC_TABLE_DATA_WIDTH)),
    758 => std_logic_vector(to_unsigned(38142, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    759 => std_logic_vector(to_unsigned(18624, LDPC_TABLE_DATA_WIDTH)),
    760 => std_logic_vector(to_unsigned(41867, LDPC_TABLE_DATA_WIDTH)),
    761 => std_logic_vector(to_unsigned(39296, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    762 => std_logic_vector(to_unsigned(37560, LDPC_TABLE_DATA_WIDTH)),
    763 => std_logic_vector(to_unsigned(14295, LDPC_TABLE_DATA_WIDTH)),
    764 => std_logic_vector(to_unsigned(16245, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    765 => std_logic_vector(to_unsigned(6821, LDPC_TABLE_DATA_WIDTH)),
    766 => std_logic_vector(to_unsigned(21679, LDPC_TABLE_DATA_WIDTH)),
    767 => std_logic_vector(to_unsigned(31570, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    768 => std_logic_vector(to_unsigned(25339, LDPC_TABLE_DATA_WIDTH)),
    769 => std_logic_vector(to_unsigned(25083, LDPC_TABLE_DATA_WIDTH)),
    770 => std_logic_vector(to_unsigned(22081, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    771 => std_logic_vector(to_unsigned(8047, LDPC_TABLE_DATA_WIDTH)),
    772 => std_logic_vector(to_unsigned(697, LDPC_TABLE_DATA_WIDTH)),
    773 => std_logic_vector(to_unsigned(35268, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    774 => std_logic_vector(to_unsigned(9884, LDPC_TABLE_DATA_WIDTH)),
    775 => std_logic_vector(to_unsigned(17073, LDPC_TABLE_DATA_WIDTH)),
    776 => std_logic_vector(to_unsigned(19995, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    777 => std_logic_vector(to_unsigned(26848, LDPC_TABLE_DATA_WIDTH)),
    778 => std_logic_vector(to_unsigned(35245, LDPC_TABLE_DATA_WIDTH)),
    779 => std_logic_vector(to_unsigned(8390, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    780 => std_logic_vector(to_unsigned(18658, LDPC_TABLE_DATA_WIDTH)),
    781 => std_logic_vector(to_unsigned(16134, LDPC_TABLE_DATA_WIDTH)),
    782 => std_logic_vector(to_unsigned(14807, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    783 => std_logic_vector(to_unsigned(12201, LDPC_TABLE_DATA_WIDTH)),
    784 => std_logic_vector(to_unsigned(32944, LDPC_TABLE_DATA_WIDTH)),
    785 => std_logic_vector(to_unsigned(5035, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    786 => std_logic_vector(to_unsigned(25236, LDPC_TABLE_DATA_WIDTH)),
    787 => std_logic_vector(to_unsigned(1216, LDPC_TABLE_DATA_WIDTH)),
    788 => std_logic_vector(to_unsigned(38986, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    789 => std_logic_vector(to_unsigned(42994, LDPC_TABLE_DATA_WIDTH)),
    790 => std_logic_vector(to_unsigned(24782, LDPC_TABLE_DATA_WIDTH)),
    791 => std_logic_vector(to_unsigned(8681, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    792 => std_logic_vector(to_unsigned(28321, LDPC_TABLE_DATA_WIDTH)),
    793 => std_logic_vector(to_unsigned(4932, LDPC_TABLE_DATA_WIDTH)),
    794 => std_logic_vector(to_unsigned(34249, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    795 => std_logic_vector(to_unsigned(4107, LDPC_TABLE_DATA_WIDTH)),
    796 => std_logic_vector(to_unsigned(29382, LDPC_TABLE_DATA_WIDTH)),
    797 => std_logic_vector(to_unsigned(32124, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    798 => std_logic_vector(to_unsigned(22157, LDPC_TABLE_DATA_WIDTH)),
    799 => std_logic_vector(to_unsigned(2624, LDPC_TABLE_DATA_WIDTH)),
    800 => std_logic_vector(to_unsigned(14468, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    801 => std_logic_vector(to_unsigned(38788, LDPC_TABLE_DATA_WIDTH)),
    802 => std_logic_vector(to_unsigned(27081, LDPC_TABLE_DATA_WIDTH)),
    803 => std_logic_vector(to_unsigned(7936, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    804 => std_logic_vector(to_unsigned(4368, LDPC_TABLE_DATA_WIDTH)),
    805 => std_logic_vector(to_unsigned(26148, LDPC_TABLE_DATA_WIDTH)),
    806 => std_logic_vector(to_unsigned(10578, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    807 => std_logic_vector(to_unsigned(25353, LDPC_TABLE_DATA_WIDTH)),
    808 => std_logic_vector(to_unsigned(4122, LDPC_TABLE_DATA_WIDTH)),
    809 => std_logic_vector(to_unsigned(39751, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C1_4
    810 => std_logic_vector(to_unsigned(23606, LDPC_TABLE_DATA_WIDTH)),
    811 => std_logic_vector(to_unsigned(36098, LDPC_TABLE_DATA_WIDTH)),
    812 => std_logic_vector(to_unsigned(1140, LDPC_TABLE_DATA_WIDTH)),
    813 => std_logic_vector(to_unsigned(28859, LDPC_TABLE_DATA_WIDTH)),
    814 => std_logic_vector(to_unsigned(18148, LDPC_TABLE_DATA_WIDTH)),
    815 => std_logic_vector(to_unsigned(18510, LDPC_TABLE_DATA_WIDTH)),
    816 => std_logic_vector(to_unsigned(6226, LDPC_TABLE_DATA_WIDTH)),
    817 => std_logic_vector(to_unsigned(540, LDPC_TABLE_DATA_WIDTH)),
    818 => std_logic_vector(to_unsigned(42014, LDPC_TABLE_DATA_WIDTH)),
    819 => std_logic_vector(to_unsigned(20879, LDPC_TABLE_DATA_WIDTH)),
    820 => std_logic_vector(to_unsigned(23802, LDPC_TABLE_DATA_WIDTH)),
    821 => std_logic_vector(to_unsigned(47088, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    822 => std_logic_vector(to_unsigned(16419, LDPC_TABLE_DATA_WIDTH)),
    823 => std_logic_vector(to_unsigned(24928, LDPC_TABLE_DATA_WIDTH)),
    824 => std_logic_vector(to_unsigned(16609, LDPC_TABLE_DATA_WIDTH)),
    825 => std_logic_vector(to_unsigned(17248, LDPC_TABLE_DATA_WIDTH)),
    826 => std_logic_vector(to_unsigned(7693, LDPC_TABLE_DATA_WIDTH)),
    827 => std_logic_vector(to_unsigned(24997, LDPC_TABLE_DATA_WIDTH)),
    828 => std_logic_vector(to_unsigned(42587, LDPC_TABLE_DATA_WIDTH)),
    829 => std_logic_vector(to_unsigned(16858, LDPC_TABLE_DATA_WIDTH)),
    830 => std_logic_vector(to_unsigned(34921, LDPC_TABLE_DATA_WIDTH)),
    831 => std_logic_vector(to_unsigned(21042, LDPC_TABLE_DATA_WIDTH)),
    832 => std_logic_vector(to_unsigned(37024, LDPC_TABLE_DATA_WIDTH)),
    833 => std_logic_vector(to_unsigned(20692, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    834 => std_logic_vector(to_unsigned(1874, LDPC_TABLE_DATA_WIDTH)),
    835 => std_logic_vector(to_unsigned(40094, LDPC_TABLE_DATA_WIDTH)),
    836 => std_logic_vector(to_unsigned(18704, LDPC_TABLE_DATA_WIDTH)),
    837 => std_logic_vector(to_unsigned(14474, LDPC_TABLE_DATA_WIDTH)),
    838 => std_logic_vector(to_unsigned(14004, LDPC_TABLE_DATA_WIDTH)),
    839 => std_logic_vector(to_unsigned(11519, LDPC_TABLE_DATA_WIDTH)),
    840 => std_logic_vector(to_unsigned(13106, LDPC_TABLE_DATA_WIDTH)),
    841 => std_logic_vector(to_unsigned(28826, LDPC_TABLE_DATA_WIDTH)),
    842 => std_logic_vector(to_unsigned(38669, LDPC_TABLE_DATA_WIDTH)),
    843 => std_logic_vector(to_unsigned(22363, LDPC_TABLE_DATA_WIDTH)),
    844 => std_logic_vector(to_unsigned(30255, LDPC_TABLE_DATA_WIDTH)),
    845 => std_logic_vector(to_unsigned(31105, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    846 => std_logic_vector(to_unsigned(22254, LDPC_TABLE_DATA_WIDTH)),
    847 => std_logic_vector(to_unsigned(40564, LDPC_TABLE_DATA_WIDTH)),
    848 => std_logic_vector(to_unsigned(22645, LDPC_TABLE_DATA_WIDTH)),
    849 => std_logic_vector(to_unsigned(22532, LDPC_TABLE_DATA_WIDTH)),
    850 => std_logic_vector(to_unsigned(6134, LDPC_TABLE_DATA_WIDTH)),
    851 => std_logic_vector(to_unsigned(9176, LDPC_TABLE_DATA_WIDTH)),
    852 => std_logic_vector(to_unsigned(39998, LDPC_TABLE_DATA_WIDTH)),
    853 => std_logic_vector(to_unsigned(23892, LDPC_TABLE_DATA_WIDTH)),
    854 => std_logic_vector(to_unsigned(8937, LDPC_TABLE_DATA_WIDTH)),
    855 => std_logic_vector(to_unsigned(15608, LDPC_TABLE_DATA_WIDTH)),
    856 => std_logic_vector(to_unsigned(16854, LDPC_TABLE_DATA_WIDTH)),
    857 => std_logic_vector(to_unsigned(31009, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    858 => std_logic_vector(to_unsigned(8037, LDPC_TABLE_DATA_WIDTH)),
    859 => std_logic_vector(to_unsigned(40401, LDPC_TABLE_DATA_WIDTH)),
    860 => std_logic_vector(to_unsigned(13550, LDPC_TABLE_DATA_WIDTH)),
    861 => std_logic_vector(to_unsigned(19526, LDPC_TABLE_DATA_WIDTH)),
    862 => std_logic_vector(to_unsigned(41902, LDPC_TABLE_DATA_WIDTH)),
    863 => std_logic_vector(to_unsigned(28782, LDPC_TABLE_DATA_WIDTH)),
    864 => std_logic_vector(to_unsigned(13304, LDPC_TABLE_DATA_WIDTH)),
    865 => std_logic_vector(to_unsigned(32796, LDPC_TABLE_DATA_WIDTH)),
    866 => std_logic_vector(to_unsigned(24679, LDPC_TABLE_DATA_WIDTH)),
    867 => std_logic_vector(to_unsigned(27140, LDPC_TABLE_DATA_WIDTH)),
    868 => std_logic_vector(to_unsigned(45980, LDPC_TABLE_DATA_WIDTH)),
    869 => std_logic_vector(to_unsigned(10021, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    870 => std_logic_vector(to_unsigned(40540, LDPC_TABLE_DATA_WIDTH)),
    871 => std_logic_vector(to_unsigned(44498, LDPC_TABLE_DATA_WIDTH)),
    872 => std_logic_vector(to_unsigned(13911, LDPC_TABLE_DATA_WIDTH)),
    873 => std_logic_vector(to_unsigned(22435, LDPC_TABLE_DATA_WIDTH)),
    874 => std_logic_vector(to_unsigned(32701, LDPC_TABLE_DATA_WIDTH)),
    875 => std_logic_vector(to_unsigned(18405, LDPC_TABLE_DATA_WIDTH)),
    876 => std_logic_vector(to_unsigned(39929, LDPC_TABLE_DATA_WIDTH)),
    877 => std_logic_vector(to_unsigned(25521, LDPC_TABLE_DATA_WIDTH)),
    878 => std_logic_vector(to_unsigned(12497, LDPC_TABLE_DATA_WIDTH)),
    879 => std_logic_vector(to_unsigned(9851, LDPC_TABLE_DATA_WIDTH)),
    880 => std_logic_vector(to_unsigned(39223, LDPC_TABLE_DATA_WIDTH)),
    881 => std_logic_vector(to_unsigned(34823, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    882 => std_logic_vector(to_unsigned(15233, LDPC_TABLE_DATA_WIDTH)),
    883 => std_logic_vector(to_unsigned(45333, LDPC_TABLE_DATA_WIDTH)),
    884 => std_logic_vector(to_unsigned(5041, LDPC_TABLE_DATA_WIDTH)),
    885 => std_logic_vector(to_unsigned(44979, LDPC_TABLE_DATA_WIDTH)),
    886 => std_logic_vector(to_unsigned(45710, LDPC_TABLE_DATA_WIDTH)),
    887 => std_logic_vector(to_unsigned(42150, LDPC_TABLE_DATA_WIDTH)),
    888 => std_logic_vector(to_unsigned(19416, LDPC_TABLE_DATA_WIDTH)),
    889 => std_logic_vector(to_unsigned(1892, LDPC_TABLE_DATA_WIDTH)),
    890 => std_logic_vector(to_unsigned(23121, LDPC_TABLE_DATA_WIDTH)),
    891 => std_logic_vector(to_unsigned(15860, LDPC_TABLE_DATA_WIDTH)),
    892 => std_logic_vector(to_unsigned(8832, LDPC_TABLE_DATA_WIDTH)),
    893 => std_logic_vector(to_unsigned(10308, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    894 => std_logic_vector(to_unsigned(10468, LDPC_TABLE_DATA_WIDTH)),
    895 => std_logic_vector(to_unsigned(44296, LDPC_TABLE_DATA_WIDTH)),
    896 => std_logic_vector(to_unsigned(3611, LDPC_TABLE_DATA_WIDTH)),
    897 => std_logic_vector(to_unsigned(1480, LDPC_TABLE_DATA_WIDTH)),
    898 => std_logic_vector(to_unsigned(37581, LDPC_TABLE_DATA_WIDTH)),
    899 => std_logic_vector(to_unsigned(32254, LDPC_TABLE_DATA_WIDTH)),
    900 => std_logic_vector(to_unsigned(13817, LDPC_TABLE_DATA_WIDTH)),
    901 => std_logic_vector(to_unsigned(6883, LDPC_TABLE_DATA_WIDTH)),
    902 => std_logic_vector(to_unsigned(32892, LDPC_TABLE_DATA_WIDTH)),
    903 => std_logic_vector(to_unsigned(40258, LDPC_TABLE_DATA_WIDTH)),
    904 => std_logic_vector(to_unsigned(46538, LDPC_TABLE_DATA_WIDTH)),
    905 => std_logic_vector(to_unsigned(11940, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    906 => std_logic_vector(to_unsigned(6705, LDPC_TABLE_DATA_WIDTH)),
    907 => std_logic_vector(to_unsigned(21634, LDPC_TABLE_DATA_WIDTH)),
    908 => std_logic_vector(to_unsigned(28150, LDPC_TABLE_DATA_WIDTH)),
    909 => std_logic_vector(to_unsigned(43757, LDPC_TABLE_DATA_WIDTH)),
    910 => std_logic_vector(to_unsigned(895, LDPC_TABLE_DATA_WIDTH)),
    911 => std_logic_vector(to_unsigned(6547, LDPC_TABLE_DATA_WIDTH)),
    912 => std_logic_vector(to_unsigned(20970, LDPC_TABLE_DATA_WIDTH)),
    913 => std_logic_vector(to_unsigned(28914, LDPC_TABLE_DATA_WIDTH)),
    914 => std_logic_vector(to_unsigned(30117, LDPC_TABLE_DATA_WIDTH)),
    915 => std_logic_vector(to_unsigned(25736, LDPC_TABLE_DATA_WIDTH)),
    916 => std_logic_vector(to_unsigned(41734, LDPC_TABLE_DATA_WIDTH)),
    917 => std_logic_vector(to_unsigned(11392, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    918 => std_logic_vector(to_unsigned(22002, LDPC_TABLE_DATA_WIDTH)),
    919 => std_logic_vector(to_unsigned(5739, LDPC_TABLE_DATA_WIDTH)),
    920 => std_logic_vector(to_unsigned(27210, LDPC_TABLE_DATA_WIDTH)),
    921 => std_logic_vector(to_unsigned(27828, LDPC_TABLE_DATA_WIDTH)),
    922 => std_logic_vector(to_unsigned(34192, LDPC_TABLE_DATA_WIDTH)),
    923 => std_logic_vector(to_unsigned(37992, LDPC_TABLE_DATA_WIDTH)),
    924 => std_logic_vector(to_unsigned(10915, LDPC_TABLE_DATA_WIDTH)),
    925 => std_logic_vector(to_unsigned(6998, LDPC_TABLE_DATA_WIDTH)),
    926 => std_logic_vector(to_unsigned(3824, LDPC_TABLE_DATA_WIDTH)),
    927 => std_logic_vector(to_unsigned(42130, LDPC_TABLE_DATA_WIDTH)),
    928 => std_logic_vector(to_unsigned(4494, LDPC_TABLE_DATA_WIDTH)),
    929 => std_logic_vector(to_unsigned(35739, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    930 => std_logic_vector(to_unsigned(8515, LDPC_TABLE_DATA_WIDTH)),
    931 => std_logic_vector(to_unsigned(1191, LDPC_TABLE_DATA_WIDTH)),
    932 => std_logic_vector(to_unsigned(13642, LDPC_TABLE_DATA_WIDTH)),
    933 => std_logic_vector(to_unsigned(30950, LDPC_TABLE_DATA_WIDTH)),
    934 => std_logic_vector(to_unsigned(25943, LDPC_TABLE_DATA_WIDTH)),
    935 => std_logic_vector(to_unsigned(12673, LDPC_TABLE_DATA_WIDTH)),
    936 => std_logic_vector(to_unsigned(16726, LDPC_TABLE_DATA_WIDTH)),
    937 => std_logic_vector(to_unsigned(34261, LDPC_TABLE_DATA_WIDTH)),
    938 => std_logic_vector(to_unsigned(31828, LDPC_TABLE_DATA_WIDTH)),
    939 => std_logic_vector(to_unsigned(3340, LDPC_TABLE_DATA_WIDTH)),
    940 => std_logic_vector(to_unsigned(8747, LDPC_TABLE_DATA_WIDTH)),
    941 => std_logic_vector(to_unsigned(39225, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    942 => std_logic_vector(to_unsigned(18979, LDPC_TABLE_DATA_WIDTH)),
    943 => std_logic_vector(to_unsigned(17058, LDPC_TABLE_DATA_WIDTH)),
    944 => std_logic_vector(to_unsigned(43130, LDPC_TABLE_DATA_WIDTH)),
    945 => std_logic_vector(to_unsigned(4246, LDPC_TABLE_DATA_WIDTH)),
    946 => std_logic_vector(to_unsigned(4793, LDPC_TABLE_DATA_WIDTH)),
    947 => std_logic_vector(to_unsigned(44030, LDPC_TABLE_DATA_WIDTH)),
    948 => std_logic_vector(to_unsigned(19454, LDPC_TABLE_DATA_WIDTH)),
    949 => std_logic_vector(to_unsigned(29511, LDPC_TABLE_DATA_WIDTH)),
    950 => std_logic_vector(to_unsigned(47929, LDPC_TABLE_DATA_WIDTH)),
    951 => std_logic_vector(to_unsigned(15174, LDPC_TABLE_DATA_WIDTH)),
    952 => std_logic_vector(to_unsigned(24333, LDPC_TABLE_DATA_WIDTH)),
    953 => std_logic_vector(to_unsigned(19354, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    954 => std_logic_vector(to_unsigned(16694, LDPC_TABLE_DATA_WIDTH)),
    955 => std_logic_vector(to_unsigned(8381, LDPC_TABLE_DATA_WIDTH)),
    956 => std_logic_vector(to_unsigned(29642, LDPC_TABLE_DATA_WIDTH)),
    957 => std_logic_vector(to_unsigned(46516, LDPC_TABLE_DATA_WIDTH)),
    958 => std_logic_vector(to_unsigned(32224, LDPC_TABLE_DATA_WIDTH)),
    959 => std_logic_vector(to_unsigned(26344, LDPC_TABLE_DATA_WIDTH)),
    960 => std_logic_vector(to_unsigned(9405, LDPC_TABLE_DATA_WIDTH)),
    961 => std_logic_vector(to_unsigned(18292, LDPC_TABLE_DATA_WIDTH)),
    962 => std_logic_vector(to_unsigned(12437, LDPC_TABLE_DATA_WIDTH)),
    963 => std_logic_vector(to_unsigned(27316, LDPC_TABLE_DATA_WIDTH)),
    964 => std_logic_vector(to_unsigned(35466, LDPC_TABLE_DATA_WIDTH)),
    965 => std_logic_vector(to_unsigned(41992, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    966 => std_logic_vector(to_unsigned(15642, LDPC_TABLE_DATA_WIDTH)),
    967 => std_logic_vector(to_unsigned(5871, LDPC_TABLE_DATA_WIDTH)),
    968 => std_logic_vector(to_unsigned(46489, LDPC_TABLE_DATA_WIDTH)),
    969 => std_logic_vector(to_unsigned(26723, LDPC_TABLE_DATA_WIDTH)),
    970 => std_logic_vector(to_unsigned(23396, LDPC_TABLE_DATA_WIDTH)),
    971 => std_logic_vector(to_unsigned(7257, LDPC_TABLE_DATA_WIDTH)),
    972 => std_logic_vector(to_unsigned(8974, LDPC_TABLE_DATA_WIDTH)),
    973 => std_logic_vector(to_unsigned(3156, LDPC_TABLE_DATA_WIDTH)),
    974 => std_logic_vector(to_unsigned(37420, LDPC_TABLE_DATA_WIDTH)),
    975 => std_logic_vector(to_unsigned(44823, LDPC_TABLE_DATA_WIDTH)),
    976 => std_logic_vector(to_unsigned(35423, LDPC_TABLE_DATA_WIDTH)),
    977 => std_logic_vector(to_unsigned(13541, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    978 => std_logic_vector(to_unsigned(42858, LDPC_TABLE_DATA_WIDTH)),
    979 => std_logic_vector(to_unsigned(32008, LDPC_TABLE_DATA_WIDTH)),
    980 => std_logic_vector(to_unsigned(41282, LDPC_TABLE_DATA_WIDTH)),
    981 => std_logic_vector(to_unsigned(38773, LDPC_TABLE_DATA_WIDTH)),
    982 => std_logic_vector(to_unsigned(26570, LDPC_TABLE_DATA_WIDTH)),
    983 => std_logic_vector(to_unsigned(2702, LDPC_TABLE_DATA_WIDTH)),
    984 => std_logic_vector(to_unsigned(27260, LDPC_TABLE_DATA_WIDTH)),
    985 => std_logic_vector(to_unsigned(46974, LDPC_TABLE_DATA_WIDTH)),
    986 => std_logic_vector(to_unsigned(1469, LDPC_TABLE_DATA_WIDTH)),
    987 => std_logic_vector(to_unsigned(20887, LDPC_TABLE_DATA_WIDTH)),
    988 => std_logic_vector(to_unsigned(27426, LDPC_TABLE_DATA_WIDTH)),
    989 => std_logic_vector(to_unsigned(38553, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    990 => std_logic_vector(to_unsigned(22152, LDPC_TABLE_DATA_WIDTH)),
    991 => std_logic_vector(to_unsigned(24261, LDPC_TABLE_DATA_WIDTH)),
    992 => std_logic_vector(to_unsigned(8297, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    993 => std_logic_vector(to_unsigned(19347, LDPC_TABLE_DATA_WIDTH)),
    994 => std_logic_vector(to_unsigned(9978, LDPC_TABLE_DATA_WIDTH)),
    995 => std_logic_vector(to_unsigned(27802, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    996 => std_logic_vector(to_unsigned(34991, LDPC_TABLE_DATA_WIDTH)),
    997 => std_logic_vector(to_unsigned(6354, LDPC_TABLE_DATA_WIDTH)),
    998 => std_logic_vector(to_unsigned(33561, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    999 => std_logic_vector(to_unsigned(29782, LDPC_TABLE_DATA_WIDTH)),
    1000 => std_logic_vector(to_unsigned(30875, LDPC_TABLE_DATA_WIDTH)),
    1001 => std_logic_vector(to_unsigned(29523, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1002 => std_logic_vector(to_unsigned(9278, LDPC_TABLE_DATA_WIDTH)),
    1003 => std_logic_vector(to_unsigned(48512, LDPC_TABLE_DATA_WIDTH)),
    1004 => std_logic_vector(to_unsigned(14349, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1005 => std_logic_vector(to_unsigned(38061, LDPC_TABLE_DATA_WIDTH)),
    1006 => std_logic_vector(to_unsigned(4165, LDPC_TABLE_DATA_WIDTH)),
    1007 => std_logic_vector(to_unsigned(43878, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1008 => std_logic_vector(to_unsigned(8548, LDPC_TABLE_DATA_WIDTH)),
    1009 => std_logic_vector(to_unsigned(33172, LDPC_TABLE_DATA_WIDTH)),
    1010 => std_logic_vector(to_unsigned(34410, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1011 => std_logic_vector(to_unsigned(22535, LDPC_TABLE_DATA_WIDTH)),
    1012 => std_logic_vector(to_unsigned(28811, LDPC_TABLE_DATA_WIDTH)),
    1013 => std_logic_vector(to_unsigned(23950, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1014 => std_logic_vector(to_unsigned(20439, LDPC_TABLE_DATA_WIDTH)),
    1015 => std_logic_vector(to_unsigned(4027, LDPC_TABLE_DATA_WIDTH)),
    1016 => std_logic_vector(to_unsigned(24186, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1017 => std_logic_vector(to_unsigned(38618, LDPC_TABLE_DATA_WIDTH)),
    1018 => std_logic_vector(to_unsigned(8187, LDPC_TABLE_DATA_WIDTH)),
    1019 => std_logic_vector(to_unsigned(30947, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1020 => std_logic_vector(to_unsigned(35538, LDPC_TABLE_DATA_WIDTH)),
    1021 => std_logic_vector(to_unsigned(43880, LDPC_TABLE_DATA_WIDTH)),
    1022 => std_logic_vector(to_unsigned(21459, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1023 => std_logic_vector(to_unsigned(7091, LDPC_TABLE_DATA_WIDTH)),
    1024 => std_logic_vector(to_unsigned(45616, LDPC_TABLE_DATA_WIDTH)),
    1025 => std_logic_vector(to_unsigned(15063, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1026 => std_logic_vector(to_unsigned(5505, LDPC_TABLE_DATA_WIDTH)),
    1027 => std_logic_vector(to_unsigned(9315, LDPC_TABLE_DATA_WIDTH)),
    1028 => std_logic_vector(to_unsigned(21908, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1029 => std_logic_vector(to_unsigned(36046, LDPC_TABLE_DATA_WIDTH)),
    1030 => std_logic_vector(to_unsigned(32914, LDPC_TABLE_DATA_WIDTH)),
    1031 => std_logic_vector(to_unsigned(11836, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1032 => std_logic_vector(to_unsigned(7304, LDPC_TABLE_DATA_WIDTH)),
    1033 => std_logic_vector(to_unsigned(39782, LDPC_TABLE_DATA_WIDTH)),
    1034 => std_logic_vector(to_unsigned(33721, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1035 => std_logic_vector(to_unsigned(16905, LDPC_TABLE_DATA_WIDTH)),
    1036 => std_logic_vector(to_unsigned(29962, LDPC_TABLE_DATA_WIDTH)),
    1037 => std_logic_vector(to_unsigned(12980, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1038 => std_logic_vector(to_unsigned(11171, LDPC_TABLE_DATA_WIDTH)),
    1039 => std_logic_vector(to_unsigned(23709, LDPC_TABLE_DATA_WIDTH)),
    1040 => std_logic_vector(to_unsigned(22460, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1041 => std_logic_vector(to_unsigned(34541, LDPC_TABLE_DATA_WIDTH)),
    1042 => std_logic_vector(to_unsigned(9937, LDPC_TABLE_DATA_WIDTH)),
    1043 => std_logic_vector(to_unsigned(44500, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1044 => std_logic_vector(to_unsigned(14035, LDPC_TABLE_DATA_WIDTH)),
    1045 => std_logic_vector(to_unsigned(47316, LDPC_TABLE_DATA_WIDTH)),
    1046 => std_logic_vector(to_unsigned(8815, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1047 => std_logic_vector(to_unsigned(15057, LDPC_TABLE_DATA_WIDTH)),
    1048 => std_logic_vector(to_unsigned(45482, LDPC_TABLE_DATA_WIDTH)),
    1049 => std_logic_vector(to_unsigned(24461, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1050 => std_logic_vector(to_unsigned(30518, LDPC_TABLE_DATA_WIDTH)),
    1051 => std_logic_vector(to_unsigned(36877, LDPC_TABLE_DATA_WIDTH)),
    1052 => std_logic_vector(to_unsigned(879, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1053 => std_logic_vector(to_unsigned(7583, LDPC_TABLE_DATA_WIDTH)),
    1054 => std_logic_vector(to_unsigned(13364, LDPC_TABLE_DATA_WIDTH)),
    1055 => std_logic_vector(to_unsigned(24332, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1056 => std_logic_vector(to_unsigned(448, LDPC_TABLE_DATA_WIDTH)),
    1057 => std_logic_vector(to_unsigned(27056, LDPC_TABLE_DATA_WIDTH)),
    1058 => std_logic_vector(to_unsigned(4682, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1059 => std_logic_vector(to_unsigned(12083, LDPC_TABLE_DATA_WIDTH)),
    1060 => std_logic_vector(to_unsigned(31378, LDPC_TABLE_DATA_WIDTH)),
    1061 => std_logic_vector(to_unsigned(21670, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1062 => std_logic_vector(to_unsigned(1159, LDPC_TABLE_DATA_WIDTH)),
    1063 => std_logic_vector(to_unsigned(18031, LDPC_TABLE_DATA_WIDTH)),
    1064 => std_logic_vector(to_unsigned(2221, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1065 => std_logic_vector(to_unsigned(17028, LDPC_TABLE_DATA_WIDTH)),
    1066 => std_logic_vector(to_unsigned(38715, LDPC_TABLE_DATA_WIDTH)),
    1067 => std_logic_vector(to_unsigned(9350, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1068 => std_logic_vector(to_unsigned(17343, LDPC_TABLE_DATA_WIDTH)),
    1069 => std_logic_vector(to_unsigned(24530, LDPC_TABLE_DATA_WIDTH)),
    1070 => std_logic_vector(to_unsigned(29574, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1071 => std_logic_vector(to_unsigned(46128, LDPC_TABLE_DATA_WIDTH)),
    1072 => std_logic_vector(to_unsigned(31039, LDPC_TABLE_DATA_WIDTH)),
    1073 => std_logic_vector(to_unsigned(32818, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1074 => std_logic_vector(to_unsigned(20373, LDPC_TABLE_DATA_WIDTH)),
    1075 => std_logic_vector(to_unsigned(36967, LDPC_TABLE_DATA_WIDTH)),
    1076 => std_logic_vector(to_unsigned(18345, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1077 => std_logic_vector(to_unsigned(46685, LDPC_TABLE_DATA_WIDTH)),
    1078 => std_logic_vector(to_unsigned(20622, LDPC_TABLE_DATA_WIDTH)),
    1079 => std_logic_vector(to_unsigned(32806, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C2_3
    1080 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    1081 => std_logic_vector(to_unsigned(10491, LDPC_TABLE_DATA_WIDTH)),
    1082 => std_logic_vector(to_unsigned(16043, LDPC_TABLE_DATA_WIDTH)),
    1083 => std_logic_vector(to_unsigned(506, LDPC_TABLE_DATA_WIDTH)),
    1084 => std_logic_vector(to_unsigned(12826, LDPC_TABLE_DATA_WIDTH)),
    1085 => std_logic_vector(to_unsigned(8065, LDPC_TABLE_DATA_WIDTH)),
    1086 => std_logic_vector(to_unsigned(8226, LDPC_TABLE_DATA_WIDTH)),
    1087 => std_logic_vector(to_unsigned(2767, LDPC_TABLE_DATA_WIDTH)),
    1088 => std_logic_vector(to_unsigned(240, LDPC_TABLE_DATA_WIDTH)),
    1089 => std_logic_vector(to_unsigned(18673, LDPC_TABLE_DATA_WIDTH)),
    1090 => std_logic_vector(to_unsigned(9279, LDPC_TABLE_DATA_WIDTH)),
    1091 => std_logic_vector(to_unsigned(10579, LDPC_TABLE_DATA_WIDTH)),
    1092 => std_logic_vector(to_unsigned(20928, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1093 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    1094 => std_logic_vector(to_unsigned(17819, LDPC_TABLE_DATA_WIDTH)),
    1095 => std_logic_vector(to_unsigned(8313, LDPC_TABLE_DATA_WIDTH)),
    1096 => std_logic_vector(to_unsigned(6433, LDPC_TABLE_DATA_WIDTH)),
    1097 => std_logic_vector(to_unsigned(6224, LDPC_TABLE_DATA_WIDTH)),
    1098 => std_logic_vector(to_unsigned(5120, LDPC_TABLE_DATA_WIDTH)),
    1099 => std_logic_vector(to_unsigned(5824, LDPC_TABLE_DATA_WIDTH)),
    1100 => std_logic_vector(to_unsigned(12812, LDPC_TABLE_DATA_WIDTH)),
    1101 => std_logic_vector(to_unsigned(17187, LDPC_TABLE_DATA_WIDTH)),
    1102 => std_logic_vector(to_unsigned(9940, LDPC_TABLE_DATA_WIDTH)),
    1103 => std_logic_vector(to_unsigned(13447, LDPC_TABLE_DATA_WIDTH)),
    1104 => std_logic_vector(to_unsigned(13825, LDPC_TABLE_DATA_WIDTH)),
    1105 => std_logic_vector(to_unsigned(18483, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1106 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    1107 => std_logic_vector(to_unsigned(17957, LDPC_TABLE_DATA_WIDTH)),
    1108 => std_logic_vector(to_unsigned(6024, LDPC_TABLE_DATA_WIDTH)),
    1109 => std_logic_vector(to_unsigned(8681, LDPC_TABLE_DATA_WIDTH)),
    1110 => std_logic_vector(to_unsigned(18628, LDPC_TABLE_DATA_WIDTH)),
    1111 => std_logic_vector(to_unsigned(12794, LDPC_TABLE_DATA_WIDTH)),
    1112 => std_logic_vector(to_unsigned(5915, LDPC_TABLE_DATA_WIDTH)),
    1113 => std_logic_vector(to_unsigned(14576, LDPC_TABLE_DATA_WIDTH)),
    1114 => std_logic_vector(to_unsigned(10970, LDPC_TABLE_DATA_WIDTH)),
    1115 => std_logic_vector(to_unsigned(12064, LDPC_TABLE_DATA_WIDTH)),
    1116 => std_logic_vector(to_unsigned(20437, LDPC_TABLE_DATA_WIDTH)),
    1117 => std_logic_vector(to_unsigned(4455, LDPC_TABLE_DATA_WIDTH)),
    1118 => std_logic_vector(to_unsigned(7151, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1119 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    1120 => std_logic_vector(to_unsigned(19777, LDPC_TABLE_DATA_WIDTH)),
    1121 => std_logic_vector(to_unsigned(6183, LDPC_TABLE_DATA_WIDTH)),
    1122 => std_logic_vector(to_unsigned(9972, LDPC_TABLE_DATA_WIDTH)),
    1123 => std_logic_vector(to_unsigned(14536, LDPC_TABLE_DATA_WIDTH)),
    1124 => std_logic_vector(to_unsigned(8182, LDPC_TABLE_DATA_WIDTH)),
    1125 => std_logic_vector(to_unsigned(17749, LDPC_TABLE_DATA_WIDTH)),
    1126 => std_logic_vector(to_unsigned(11341, LDPC_TABLE_DATA_WIDTH)),
    1127 => std_logic_vector(to_unsigned(5556, LDPC_TABLE_DATA_WIDTH)),
    1128 => std_logic_vector(to_unsigned(4379, LDPC_TABLE_DATA_WIDTH)),
    1129 => std_logic_vector(to_unsigned(17434, LDPC_TABLE_DATA_WIDTH)),
    1130 => std_logic_vector(to_unsigned(15477, LDPC_TABLE_DATA_WIDTH)),
    1131 => std_logic_vector(to_unsigned(18532, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1132 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    1133 => std_logic_vector(to_unsigned(4651, LDPC_TABLE_DATA_WIDTH)),
    1134 => std_logic_vector(to_unsigned(19689, LDPC_TABLE_DATA_WIDTH)),
    1135 => std_logic_vector(to_unsigned(1608, LDPC_TABLE_DATA_WIDTH)),
    1136 => std_logic_vector(to_unsigned(659, LDPC_TABLE_DATA_WIDTH)),
    1137 => std_logic_vector(to_unsigned(16707, LDPC_TABLE_DATA_WIDTH)),
    1138 => std_logic_vector(to_unsigned(14335, LDPC_TABLE_DATA_WIDTH)),
    1139 => std_logic_vector(to_unsigned(6143, LDPC_TABLE_DATA_WIDTH)),
    1140 => std_logic_vector(to_unsigned(3058, LDPC_TABLE_DATA_WIDTH)),
    1141 => std_logic_vector(to_unsigned(14618, LDPC_TABLE_DATA_WIDTH)),
    1142 => std_logic_vector(to_unsigned(17894, LDPC_TABLE_DATA_WIDTH)),
    1143 => std_logic_vector(to_unsigned(20684, LDPC_TABLE_DATA_WIDTH)),
    1144 => std_logic_vector(to_unsigned(5306, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1145 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    1146 => std_logic_vector(to_unsigned(9778, LDPC_TABLE_DATA_WIDTH)),
    1147 => std_logic_vector(to_unsigned(2552, LDPC_TABLE_DATA_WIDTH)),
    1148 => std_logic_vector(to_unsigned(12096, LDPC_TABLE_DATA_WIDTH)),
    1149 => std_logic_vector(to_unsigned(12369, LDPC_TABLE_DATA_WIDTH)),
    1150 => std_logic_vector(to_unsigned(15198, LDPC_TABLE_DATA_WIDTH)),
    1151 => std_logic_vector(to_unsigned(16890, LDPC_TABLE_DATA_WIDTH)),
    1152 => std_logic_vector(to_unsigned(4851, LDPC_TABLE_DATA_WIDTH)),
    1153 => std_logic_vector(to_unsigned(3109, LDPC_TABLE_DATA_WIDTH)),
    1154 => std_logic_vector(to_unsigned(1700, LDPC_TABLE_DATA_WIDTH)),
    1155 => std_logic_vector(to_unsigned(18725, LDPC_TABLE_DATA_WIDTH)),
    1156 => std_logic_vector(to_unsigned(1997, LDPC_TABLE_DATA_WIDTH)),
    1157 => std_logic_vector(to_unsigned(15882, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1158 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    1159 => std_logic_vector(to_unsigned(486, LDPC_TABLE_DATA_WIDTH)),
    1160 => std_logic_vector(to_unsigned(6111, LDPC_TABLE_DATA_WIDTH)),
    1161 => std_logic_vector(to_unsigned(13743, LDPC_TABLE_DATA_WIDTH)),
    1162 => std_logic_vector(to_unsigned(11537, LDPC_TABLE_DATA_WIDTH)),
    1163 => std_logic_vector(to_unsigned(5591, LDPC_TABLE_DATA_WIDTH)),
    1164 => std_logic_vector(to_unsigned(7433, LDPC_TABLE_DATA_WIDTH)),
    1165 => std_logic_vector(to_unsigned(15227, LDPC_TABLE_DATA_WIDTH)),
    1166 => std_logic_vector(to_unsigned(14145, LDPC_TABLE_DATA_WIDTH)),
    1167 => std_logic_vector(to_unsigned(1483, LDPC_TABLE_DATA_WIDTH)),
    1168 => std_logic_vector(to_unsigned(3887, LDPC_TABLE_DATA_WIDTH)),
    1169 => std_logic_vector(to_unsigned(17431, LDPC_TABLE_DATA_WIDTH)),
    1170 => std_logic_vector(to_unsigned(12430, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1171 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    1172 => std_logic_vector(to_unsigned(20647, LDPC_TABLE_DATA_WIDTH)),
    1173 => std_logic_vector(to_unsigned(14311, LDPC_TABLE_DATA_WIDTH)),
    1174 => std_logic_vector(to_unsigned(11734, LDPC_TABLE_DATA_WIDTH)),
    1175 => std_logic_vector(to_unsigned(4180, LDPC_TABLE_DATA_WIDTH)),
    1176 => std_logic_vector(to_unsigned(8110, LDPC_TABLE_DATA_WIDTH)),
    1177 => std_logic_vector(to_unsigned(5525, LDPC_TABLE_DATA_WIDTH)),
    1178 => std_logic_vector(to_unsigned(12141, LDPC_TABLE_DATA_WIDTH)),
    1179 => std_logic_vector(to_unsigned(15761, LDPC_TABLE_DATA_WIDTH)),
    1180 => std_logic_vector(to_unsigned(18661, LDPC_TABLE_DATA_WIDTH)),
    1181 => std_logic_vector(to_unsigned(18441, LDPC_TABLE_DATA_WIDTH)),
    1182 => std_logic_vector(to_unsigned(10569, LDPC_TABLE_DATA_WIDTH)),
    1183 => std_logic_vector(to_unsigned(8192, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1184 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    1185 => std_logic_vector(to_unsigned(3791, LDPC_TABLE_DATA_WIDTH)),
    1186 => std_logic_vector(to_unsigned(14759, LDPC_TABLE_DATA_WIDTH)),
    1187 => std_logic_vector(to_unsigned(15264, LDPC_TABLE_DATA_WIDTH)),
    1188 => std_logic_vector(to_unsigned(19918, LDPC_TABLE_DATA_WIDTH)),
    1189 => std_logic_vector(to_unsigned(10132, LDPC_TABLE_DATA_WIDTH)),
    1190 => std_logic_vector(to_unsigned(9062, LDPC_TABLE_DATA_WIDTH)),
    1191 => std_logic_vector(to_unsigned(10010, LDPC_TABLE_DATA_WIDTH)),
    1192 => std_logic_vector(to_unsigned(12786, LDPC_TABLE_DATA_WIDTH)),
    1193 => std_logic_vector(to_unsigned(10675, LDPC_TABLE_DATA_WIDTH)),
    1194 => std_logic_vector(to_unsigned(9682, LDPC_TABLE_DATA_WIDTH)),
    1195 => std_logic_vector(to_unsigned(19246, LDPC_TABLE_DATA_WIDTH)),
    1196 => std_logic_vector(to_unsigned(5454, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1197 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    1198 => std_logic_vector(to_unsigned(19525, LDPC_TABLE_DATA_WIDTH)),
    1199 => std_logic_vector(to_unsigned(9485, LDPC_TABLE_DATA_WIDTH)),
    1200 => std_logic_vector(to_unsigned(7777, LDPC_TABLE_DATA_WIDTH)),
    1201 => std_logic_vector(to_unsigned(19999, LDPC_TABLE_DATA_WIDTH)),
    1202 => std_logic_vector(to_unsigned(8378, LDPC_TABLE_DATA_WIDTH)),
    1203 => std_logic_vector(to_unsigned(9209, LDPC_TABLE_DATA_WIDTH)),
    1204 => std_logic_vector(to_unsigned(3163, LDPC_TABLE_DATA_WIDTH)),
    1205 => std_logic_vector(to_unsigned(20232, LDPC_TABLE_DATA_WIDTH)),
    1206 => std_logic_vector(to_unsigned(6690, LDPC_TABLE_DATA_WIDTH)),
    1207 => std_logic_vector(to_unsigned(16518, LDPC_TABLE_DATA_WIDTH)),
    1208 => std_logic_vector(to_unsigned(716, LDPC_TABLE_DATA_WIDTH)),
    1209 => std_logic_vector(to_unsigned(7353, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1210 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    1211 => std_logic_vector(to_unsigned(4588, LDPC_TABLE_DATA_WIDTH)),
    1212 => std_logic_vector(to_unsigned(6709, LDPC_TABLE_DATA_WIDTH)),
    1213 => std_logic_vector(to_unsigned(20202, LDPC_TABLE_DATA_WIDTH)),
    1214 => std_logic_vector(to_unsigned(10905, LDPC_TABLE_DATA_WIDTH)),
    1215 => std_logic_vector(to_unsigned(915, LDPC_TABLE_DATA_WIDTH)),
    1216 => std_logic_vector(to_unsigned(4317, LDPC_TABLE_DATA_WIDTH)),
    1217 => std_logic_vector(to_unsigned(11073, LDPC_TABLE_DATA_WIDTH)),
    1218 => std_logic_vector(to_unsigned(13576, LDPC_TABLE_DATA_WIDTH)),
    1219 => std_logic_vector(to_unsigned(16433, LDPC_TABLE_DATA_WIDTH)),
    1220 => std_logic_vector(to_unsigned(368, LDPC_TABLE_DATA_WIDTH)),
    1221 => std_logic_vector(to_unsigned(3508, LDPC_TABLE_DATA_WIDTH)),
    1222 => std_logic_vector(to_unsigned(21171, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1223 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    1224 => std_logic_vector(to_unsigned(14072, LDPC_TABLE_DATA_WIDTH)),
    1225 => std_logic_vector(to_unsigned(4033, LDPC_TABLE_DATA_WIDTH)),
    1226 => std_logic_vector(to_unsigned(19959, LDPC_TABLE_DATA_WIDTH)),
    1227 => std_logic_vector(to_unsigned(12608, LDPC_TABLE_DATA_WIDTH)),
    1228 => std_logic_vector(to_unsigned(631, LDPC_TABLE_DATA_WIDTH)),
    1229 => std_logic_vector(to_unsigned(19494, LDPC_TABLE_DATA_WIDTH)),
    1230 => std_logic_vector(to_unsigned(14160, LDPC_TABLE_DATA_WIDTH)),
    1231 => std_logic_vector(to_unsigned(8249, LDPC_TABLE_DATA_WIDTH)),
    1232 => std_logic_vector(to_unsigned(10223, LDPC_TABLE_DATA_WIDTH)),
    1233 => std_logic_vector(to_unsigned(21504, LDPC_TABLE_DATA_WIDTH)),
    1234 => std_logic_vector(to_unsigned(12395, LDPC_TABLE_DATA_WIDTH)),
    1235 => std_logic_vector(to_unsigned(4322, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1236 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    1237 => std_logic_vector(to_unsigned(13800, LDPC_TABLE_DATA_WIDTH)),
    1238 => std_logic_vector(to_unsigned(14161, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1239 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    1240 => std_logic_vector(to_unsigned(2948, LDPC_TABLE_DATA_WIDTH)),
    1241 => std_logic_vector(to_unsigned(9647, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1242 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    1243 => std_logic_vector(to_unsigned(14693, LDPC_TABLE_DATA_WIDTH)),
    1244 => std_logic_vector(to_unsigned(16027, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1245 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    1246 => std_logic_vector(to_unsigned(20506, LDPC_TABLE_DATA_WIDTH)),
    1247 => std_logic_vector(to_unsigned(11082, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1248 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    1249 => std_logic_vector(to_unsigned(1143, LDPC_TABLE_DATA_WIDTH)),
    1250 => std_logic_vector(to_unsigned(9020, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1251 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    1252 => std_logic_vector(to_unsigned(13501, LDPC_TABLE_DATA_WIDTH)),
    1253 => std_logic_vector(to_unsigned(4014, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1254 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    1255 => std_logic_vector(to_unsigned(1548, LDPC_TABLE_DATA_WIDTH)),
    1256 => std_logic_vector(to_unsigned(2190, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1257 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    1258 => std_logic_vector(to_unsigned(12216, LDPC_TABLE_DATA_WIDTH)),
    1259 => std_logic_vector(to_unsigned(21556, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1260 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    1261 => std_logic_vector(to_unsigned(2095, LDPC_TABLE_DATA_WIDTH)),
    1262 => std_logic_vector(to_unsigned(19897, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1263 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    1264 => std_logic_vector(to_unsigned(4189, LDPC_TABLE_DATA_WIDTH)),
    1265 => std_logic_vector(to_unsigned(7958, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1266 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    1267 => std_logic_vector(to_unsigned(15940, LDPC_TABLE_DATA_WIDTH)),
    1268 => std_logic_vector(to_unsigned(10048, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1269 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    1270 => std_logic_vector(to_unsigned(515, LDPC_TABLE_DATA_WIDTH)),
    1271 => std_logic_vector(to_unsigned(12614, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1272 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    1273 => std_logic_vector(to_unsigned(8501, LDPC_TABLE_DATA_WIDTH)),
    1274 => std_logic_vector(to_unsigned(8450, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1275 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    1276 => std_logic_vector(to_unsigned(17595, LDPC_TABLE_DATA_WIDTH)),
    1277 => std_logic_vector(to_unsigned(16784, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1278 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    1279 => std_logic_vector(to_unsigned(5913, LDPC_TABLE_DATA_WIDTH)),
    1280 => std_logic_vector(to_unsigned(8495, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1281 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    1282 => std_logic_vector(to_unsigned(16394, LDPC_TABLE_DATA_WIDTH)),
    1283 => std_logic_vector(to_unsigned(10423, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1284 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    1285 => std_logic_vector(to_unsigned(7409, LDPC_TABLE_DATA_WIDTH)),
    1286 => std_logic_vector(to_unsigned(6981, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1287 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    1288 => std_logic_vector(to_unsigned(6678, LDPC_TABLE_DATA_WIDTH)),
    1289 => std_logic_vector(to_unsigned(15939, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1290 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    1291 => std_logic_vector(to_unsigned(20344, LDPC_TABLE_DATA_WIDTH)),
    1292 => std_logic_vector(to_unsigned(12987, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1293 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    1294 => std_logic_vector(to_unsigned(2510, LDPC_TABLE_DATA_WIDTH)),
    1295 => std_logic_vector(to_unsigned(14588, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1296 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    1297 => std_logic_vector(to_unsigned(17918, LDPC_TABLE_DATA_WIDTH)),
    1298 => std_logic_vector(to_unsigned(6655, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1299 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    1300 => std_logic_vector(to_unsigned(6703, LDPC_TABLE_DATA_WIDTH)),
    1301 => std_logic_vector(to_unsigned(19451, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1302 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    1303 => std_logic_vector(to_unsigned(496, LDPC_TABLE_DATA_WIDTH)),
    1304 => std_logic_vector(to_unsigned(4217, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1305 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    1306 => std_logic_vector(to_unsigned(7290, LDPC_TABLE_DATA_WIDTH)),
    1307 => std_logic_vector(to_unsigned(5766, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1308 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    1309 => std_logic_vector(to_unsigned(10521, LDPC_TABLE_DATA_WIDTH)),
    1310 => std_logic_vector(to_unsigned(8925, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1311 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    1312 => std_logic_vector(to_unsigned(20379, LDPC_TABLE_DATA_WIDTH)),
    1313 => std_logic_vector(to_unsigned(11905, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1314 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    1315 => std_logic_vector(to_unsigned(4090, LDPC_TABLE_DATA_WIDTH)),
    1316 => std_logic_vector(to_unsigned(5838, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1317 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    1318 => std_logic_vector(to_unsigned(19082, LDPC_TABLE_DATA_WIDTH)),
    1319 => std_logic_vector(to_unsigned(17040, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1320 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    1321 => std_logic_vector(to_unsigned(20233, LDPC_TABLE_DATA_WIDTH)),
    1322 => std_logic_vector(to_unsigned(12352, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1323 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    1324 => std_logic_vector(to_unsigned(19365, LDPC_TABLE_DATA_WIDTH)),
    1325 => std_logic_vector(to_unsigned(19546, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1326 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    1327 => std_logic_vector(to_unsigned(6249, LDPC_TABLE_DATA_WIDTH)),
    1328 => std_logic_vector(to_unsigned(19030, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1329 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    1330 => std_logic_vector(to_unsigned(11037, LDPC_TABLE_DATA_WIDTH)),
    1331 => std_logic_vector(to_unsigned(19193, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1332 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    1333 => std_logic_vector(to_unsigned(19760, LDPC_TABLE_DATA_WIDTH)),
    1334 => std_logic_vector(to_unsigned(11772, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1335 => std_logic_vector(to_unsigned(45, LDPC_TABLE_DATA_WIDTH)),
    1336 => std_logic_vector(to_unsigned(19644, LDPC_TABLE_DATA_WIDTH)),
    1337 => std_logic_vector(to_unsigned(7428, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1338 => std_logic_vector(to_unsigned(46, LDPC_TABLE_DATA_WIDTH)),
    1339 => std_logic_vector(to_unsigned(16076, LDPC_TABLE_DATA_WIDTH)),
    1340 => std_logic_vector(to_unsigned(3521, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1341 => std_logic_vector(to_unsigned(47, LDPC_TABLE_DATA_WIDTH)),
    1342 => std_logic_vector(to_unsigned(11779, LDPC_TABLE_DATA_WIDTH)),
    1343 => std_logic_vector(to_unsigned(21062, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1344 => std_logic_vector(to_unsigned(48, LDPC_TABLE_DATA_WIDTH)),
    1345 => std_logic_vector(to_unsigned(13062, LDPC_TABLE_DATA_WIDTH)),
    1346 => std_logic_vector(to_unsigned(9682, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1347 => std_logic_vector(to_unsigned(49, LDPC_TABLE_DATA_WIDTH)),
    1348 => std_logic_vector(to_unsigned(8934, LDPC_TABLE_DATA_WIDTH)),
    1349 => std_logic_vector(to_unsigned(5217, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1350 => std_logic_vector(to_unsigned(50, LDPC_TABLE_DATA_WIDTH)),
    1351 => std_logic_vector(to_unsigned(11087, LDPC_TABLE_DATA_WIDTH)),
    1352 => std_logic_vector(to_unsigned(3319, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1353 => std_logic_vector(to_unsigned(51, LDPC_TABLE_DATA_WIDTH)),
    1354 => std_logic_vector(to_unsigned(18892, LDPC_TABLE_DATA_WIDTH)),
    1355 => std_logic_vector(to_unsigned(4356, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1356 => std_logic_vector(to_unsigned(52, LDPC_TABLE_DATA_WIDTH)),
    1357 => std_logic_vector(to_unsigned(7894, LDPC_TABLE_DATA_WIDTH)),
    1358 => std_logic_vector(to_unsigned(3898, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1359 => std_logic_vector(to_unsigned(53, LDPC_TABLE_DATA_WIDTH)),
    1360 => std_logic_vector(to_unsigned(5963, LDPC_TABLE_DATA_WIDTH)),
    1361 => std_logic_vector(to_unsigned(4360, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1362 => std_logic_vector(to_unsigned(54, LDPC_TABLE_DATA_WIDTH)),
    1363 => std_logic_vector(to_unsigned(7346, LDPC_TABLE_DATA_WIDTH)),
    1364 => std_logic_vector(to_unsigned(11726, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1365 => std_logic_vector(to_unsigned(55, LDPC_TABLE_DATA_WIDTH)),
    1366 => std_logic_vector(to_unsigned(5182, LDPC_TABLE_DATA_WIDTH)),
    1367 => std_logic_vector(to_unsigned(5609, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1368 => std_logic_vector(to_unsigned(56, LDPC_TABLE_DATA_WIDTH)),
    1369 => std_logic_vector(to_unsigned(2412, LDPC_TABLE_DATA_WIDTH)),
    1370 => std_logic_vector(to_unsigned(17295, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1371 => std_logic_vector(to_unsigned(57, LDPC_TABLE_DATA_WIDTH)),
    1372 => std_logic_vector(to_unsigned(9845, LDPC_TABLE_DATA_WIDTH)),
    1373 => std_logic_vector(to_unsigned(20494, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1374 => std_logic_vector(to_unsigned(58, LDPC_TABLE_DATA_WIDTH)),
    1375 => std_logic_vector(to_unsigned(6687, LDPC_TABLE_DATA_WIDTH)),
    1376 => std_logic_vector(to_unsigned(1864, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1377 => std_logic_vector(to_unsigned(59, LDPC_TABLE_DATA_WIDTH)),
    1378 => std_logic_vector(to_unsigned(20564, LDPC_TABLE_DATA_WIDTH)),
    1379 => std_logic_vector(to_unsigned(5216, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1380 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    1381 => std_logic_vector(to_unsigned(18226, LDPC_TABLE_DATA_WIDTH)),
    1382 => std_logic_vector(to_unsigned(17207, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1383 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    1384 => std_logic_vector(to_unsigned(9380, LDPC_TABLE_DATA_WIDTH)),
    1385 => std_logic_vector(to_unsigned(8266, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1386 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    1387 => std_logic_vector(to_unsigned(7073, LDPC_TABLE_DATA_WIDTH)),
    1388 => std_logic_vector(to_unsigned(3065, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1389 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    1390 => std_logic_vector(to_unsigned(18252, LDPC_TABLE_DATA_WIDTH)),
    1391 => std_logic_vector(to_unsigned(13437, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1392 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    1393 => std_logic_vector(to_unsigned(9161, LDPC_TABLE_DATA_WIDTH)),
    1394 => std_logic_vector(to_unsigned(15642, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1395 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    1396 => std_logic_vector(to_unsigned(10714, LDPC_TABLE_DATA_WIDTH)),
    1397 => std_logic_vector(to_unsigned(10153, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1398 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    1399 => std_logic_vector(to_unsigned(11585, LDPC_TABLE_DATA_WIDTH)),
    1400 => std_logic_vector(to_unsigned(9078, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1401 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    1402 => std_logic_vector(to_unsigned(5359, LDPC_TABLE_DATA_WIDTH)),
    1403 => std_logic_vector(to_unsigned(9418, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1404 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    1405 => std_logic_vector(to_unsigned(9024, LDPC_TABLE_DATA_WIDTH)),
    1406 => std_logic_vector(to_unsigned(9515, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1407 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    1408 => std_logic_vector(to_unsigned(1206, LDPC_TABLE_DATA_WIDTH)),
    1409 => std_logic_vector(to_unsigned(16354, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1410 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    1411 => std_logic_vector(to_unsigned(14994, LDPC_TABLE_DATA_WIDTH)),
    1412 => std_logic_vector(to_unsigned(1102, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1413 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    1414 => std_logic_vector(to_unsigned(9375, LDPC_TABLE_DATA_WIDTH)),
    1415 => std_logic_vector(to_unsigned(20796, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1416 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    1417 => std_logic_vector(to_unsigned(15964, LDPC_TABLE_DATA_WIDTH)),
    1418 => std_logic_vector(to_unsigned(6027, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1419 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    1420 => std_logic_vector(to_unsigned(14789, LDPC_TABLE_DATA_WIDTH)),
    1421 => std_logic_vector(to_unsigned(6452, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1422 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    1423 => std_logic_vector(to_unsigned(8002, LDPC_TABLE_DATA_WIDTH)),
    1424 => std_logic_vector(to_unsigned(18591, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1425 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    1426 => std_logic_vector(to_unsigned(14742, LDPC_TABLE_DATA_WIDTH)),
    1427 => std_logic_vector(to_unsigned(14089, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1428 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    1429 => std_logic_vector(to_unsigned(253, LDPC_TABLE_DATA_WIDTH)),
    1430 => std_logic_vector(to_unsigned(3045, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1431 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    1432 => std_logic_vector(to_unsigned(1274, LDPC_TABLE_DATA_WIDTH)),
    1433 => std_logic_vector(to_unsigned(19286, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1434 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    1435 => std_logic_vector(to_unsigned(14777, LDPC_TABLE_DATA_WIDTH)),
    1436 => std_logic_vector(to_unsigned(2044, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1437 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    1438 => std_logic_vector(to_unsigned(13920, LDPC_TABLE_DATA_WIDTH)),
    1439 => std_logic_vector(to_unsigned(9900, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1440 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    1441 => std_logic_vector(to_unsigned(452, LDPC_TABLE_DATA_WIDTH)),
    1442 => std_logic_vector(to_unsigned(7374, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1443 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    1444 => std_logic_vector(to_unsigned(18206, LDPC_TABLE_DATA_WIDTH)),
    1445 => std_logic_vector(to_unsigned(9921, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1446 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    1447 => std_logic_vector(to_unsigned(6131, LDPC_TABLE_DATA_WIDTH)),
    1448 => std_logic_vector(to_unsigned(5414, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1449 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    1450 => std_logic_vector(to_unsigned(10077, LDPC_TABLE_DATA_WIDTH)),
    1451 => std_logic_vector(to_unsigned(9726, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1452 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    1453 => std_logic_vector(to_unsigned(12045, LDPC_TABLE_DATA_WIDTH)),
    1454 => std_logic_vector(to_unsigned(5479, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1455 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    1456 => std_logic_vector(to_unsigned(4322, LDPC_TABLE_DATA_WIDTH)),
    1457 => std_logic_vector(to_unsigned(7990, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1458 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    1459 => std_logic_vector(to_unsigned(15616, LDPC_TABLE_DATA_WIDTH)),
    1460 => std_logic_vector(to_unsigned(5550, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1461 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    1462 => std_logic_vector(to_unsigned(15561, LDPC_TABLE_DATA_WIDTH)),
    1463 => std_logic_vector(to_unsigned(10661, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1464 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    1465 => std_logic_vector(to_unsigned(20718, LDPC_TABLE_DATA_WIDTH)),
    1466 => std_logic_vector(to_unsigned(7387, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1467 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    1468 => std_logic_vector(to_unsigned(2518, LDPC_TABLE_DATA_WIDTH)),
    1469 => std_logic_vector(to_unsigned(18804, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1470 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    1471 => std_logic_vector(to_unsigned(8984, LDPC_TABLE_DATA_WIDTH)),
    1472 => std_logic_vector(to_unsigned(2600, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1473 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    1474 => std_logic_vector(to_unsigned(6516, LDPC_TABLE_DATA_WIDTH)),
    1475 => std_logic_vector(to_unsigned(17909, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1476 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    1477 => std_logic_vector(to_unsigned(11148, LDPC_TABLE_DATA_WIDTH)),
    1478 => std_logic_vector(to_unsigned(98, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1479 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    1480 => std_logic_vector(to_unsigned(20559, LDPC_TABLE_DATA_WIDTH)),
    1481 => std_logic_vector(to_unsigned(3704, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1482 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    1483 => std_logic_vector(to_unsigned(7510, LDPC_TABLE_DATA_WIDTH)),
    1484 => std_logic_vector(to_unsigned(1569, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1485 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    1486 => std_logic_vector(to_unsigned(16000, LDPC_TABLE_DATA_WIDTH)),
    1487 => std_logic_vector(to_unsigned(11692, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1488 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    1489 => std_logic_vector(to_unsigned(9147, LDPC_TABLE_DATA_WIDTH)),
    1490 => std_logic_vector(to_unsigned(10303, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1491 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    1492 => std_logic_vector(to_unsigned(16650, LDPC_TABLE_DATA_WIDTH)),
    1493 => std_logic_vector(to_unsigned(191, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1494 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    1495 => std_logic_vector(to_unsigned(15577, LDPC_TABLE_DATA_WIDTH)),
    1496 => std_logic_vector(to_unsigned(18685, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1497 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    1498 => std_logic_vector(to_unsigned(17167, LDPC_TABLE_DATA_WIDTH)),
    1499 => std_logic_vector(to_unsigned(20917, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1500 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    1501 => std_logic_vector(to_unsigned(4256, LDPC_TABLE_DATA_WIDTH)),
    1502 => std_logic_vector(to_unsigned(3391, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1503 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    1504 => std_logic_vector(to_unsigned(20092, LDPC_TABLE_DATA_WIDTH)),
    1505 => std_logic_vector(to_unsigned(17219, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1506 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    1507 => std_logic_vector(to_unsigned(9218, LDPC_TABLE_DATA_WIDTH)),
    1508 => std_logic_vector(to_unsigned(5056, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1509 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    1510 => std_logic_vector(to_unsigned(18429, LDPC_TABLE_DATA_WIDTH)),
    1511 => std_logic_vector(to_unsigned(8472, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1512 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    1513 => std_logic_vector(to_unsigned(12093, LDPC_TABLE_DATA_WIDTH)),
    1514 => std_logic_vector(to_unsigned(20753, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1515 => std_logic_vector(to_unsigned(45, LDPC_TABLE_DATA_WIDTH)),
    1516 => std_logic_vector(to_unsigned(16345, LDPC_TABLE_DATA_WIDTH)),
    1517 => std_logic_vector(to_unsigned(12748, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1518 => std_logic_vector(to_unsigned(46, LDPC_TABLE_DATA_WIDTH)),
    1519 => std_logic_vector(to_unsigned(16023, LDPC_TABLE_DATA_WIDTH)),
    1520 => std_logic_vector(to_unsigned(11095, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1521 => std_logic_vector(to_unsigned(47, LDPC_TABLE_DATA_WIDTH)),
    1522 => std_logic_vector(to_unsigned(5048, LDPC_TABLE_DATA_WIDTH)),
    1523 => std_logic_vector(to_unsigned(17595, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1524 => std_logic_vector(to_unsigned(48, LDPC_TABLE_DATA_WIDTH)),
    1525 => std_logic_vector(to_unsigned(18995, LDPC_TABLE_DATA_WIDTH)),
    1526 => std_logic_vector(to_unsigned(4817, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1527 => std_logic_vector(to_unsigned(49, LDPC_TABLE_DATA_WIDTH)),
    1528 => std_logic_vector(to_unsigned(16483, LDPC_TABLE_DATA_WIDTH)),
    1529 => std_logic_vector(to_unsigned(3536, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1530 => std_logic_vector(to_unsigned(50, LDPC_TABLE_DATA_WIDTH)),
    1531 => std_logic_vector(to_unsigned(1439, LDPC_TABLE_DATA_WIDTH)),
    1532 => std_logic_vector(to_unsigned(16148, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1533 => std_logic_vector(to_unsigned(51, LDPC_TABLE_DATA_WIDTH)),
    1534 => std_logic_vector(to_unsigned(3661, LDPC_TABLE_DATA_WIDTH)),
    1535 => std_logic_vector(to_unsigned(3039, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1536 => std_logic_vector(to_unsigned(52, LDPC_TABLE_DATA_WIDTH)),
    1537 => std_logic_vector(to_unsigned(19010, LDPC_TABLE_DATA_WIDTH)),
    1538 => std_logic_vector(to_unsigned(18121, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1539 => std_logic_vector(to_unsigned(53, LDPC_TABLE_DATA_WIDTH)),
    1540 => std_logic_vector(to_unsigned(8968, LDPC_TABLE_DATA_WIDTH)),
    1541 => std_logic_vector(to_unsigned(11793, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1542 => std_logic_vector(to_unsigned(54, LDPC_TABLE_DATA_WIDTH)),
    1543 => std_logic_vector(to_unsigned(13427, LDPC_TABLE_DATA_WIDTH)),
    1544 => std_logic_vector(to_unsigned(18003, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1545 => std_logic_vector(to_unsigned(55, LDPC_TABLE_DATA_WIDTH)),
    1546 => std_logic_vector(to_unsigned(5303, LDPC_TABLE_DATA_WIDTH)),
    1547 => std_logic_vector(to_unsigned(3083, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1548 => std_logic_vector(to_unsigned(56, LDPC_TABLE_DATA_WIDTH)),
    1549 => std_logic_vector(to_unsigned(531, LDPC_TABLE_DATA_WIDTH)),
    1550 => std_logic_vector(to_unsigned(16668, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1551 => std_logic_vector(to_unsigned(57, LDPC_TABLE_DATA_WIDTH)),
    1552 => std_logic_vector(to_unsigned(4771, LDPC_TABLE_DATA_WIDTH)),
    1553 => std_logic_vector(to_unsigned(6722, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1554 => std_logic_vector(to_unsigned(58, LDPC_TABLE_DATA_WIDTH)),
    1555 => std_logic_vector(to_unsigned(5695, LDPC_TABLE_DATA_WIDTH)),
    1556 => std_logic_vector(to_unsigned(7960, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1557 => std_logic_vector(to_unsigned(59, LDPC_TABLE_DATA_WIDTH)),
    1558 => std_logic_vector(to_unsigned(3589, LDPC_TABLE_DATA_WIDTH)),
    1559 => std_logic_vector(to_unsigned(14630, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C2_5
    1560 => std_logic_vector(to_unsigned(31413, LDPC_TABLE_DATA_WIDTH)),
    1561 => std_logic_vector(to_unsigned(18834, LDPC_TABLE_DATA_WIDTH)),
    1562 => std_logic_vector(to_unsigned(28884, LDPC_TABLE_DATA_WIDTH)),
    1563 => std_logic_vector(to_unsigned(947, LDPC_TABLE_DATA_WIDTH)),
    1564 => std_logic_vector(to_unsigned(23050, LDPC_TABLE_DATA_WIDTH)),
    1565 => std_logic_vector(to_unsigned(14484, LDPC_TABLE_DATA_WIDTH)),
    1566 => std_logic_vector(to_unsigned(14809, LDPC_TABLE_DATA_WIDTH)),
    1567 => std_logic_vector(to_unsigned(4968, LDPC_TABLE_DATA_WIDTH)),
    1568 => std_logic_vector(to_unsigned(455, LDPC_TABLE_DATA_WIDTH)),
    1569 => std_logic_vector(to_unsigned(33659, LDPC_TABLE_DATA_WIDTH)),
    1570 => std_logic_vector(to_unsigned(16666, LDPC_TABLE_DATA_WIDTH)),
    1571 => std_logic_vector(to_unsigned(19008, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1572 => std_logic_vector(to_unsigned(13172, LDPC_TABLE_DATA_WIDTH)),
    1573 => std_logic_vector(to_unsigned(19939, LDPC_TABLE_DATA_WIDTH)),
    1574 => std_logic_vector(to_unsigned(13354, LDPC_TABLE_DATA_WIDTH)),
    1575 => std_logic_vector(to_unsigned(13719, LDPC_TABLE_DATA_WIDTH)),
    1576 => std_logic_vector(to_unsigned(6132, LDPC_TABLE_DATA_WIDTH)),
    1577 => std_logic_vector(to_unsigned(20086, LDPC_TABLE_DATA_WIDTH)),
    1578 => std_logic_vector(to_unsigned(34040, LDPC_TABLE_DATA_WIDTH)),
    1579 => std_logic_vector(to_unsigned(13442, LDPC_TABLE_DATA_WIDTH)),
    1580 => std_logic_vector(to_unsigned(27958, LDPC_TABLE_DATA_WIDTH)),
    1581 => std_logic_vector(to_unsigned(16813, LDPC_TABLE_DATA_WIDTH)),
    1582 => std_logic_vector(to_unsigned(29619, LDPC_TABLE_DATA_WIDTH)),
    1583 => std_logic_vector(to_unsigned(16553, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1584 => std_logic_vector(to_unsigned(1499, LDPC_TABLE_DATA_WIDTH)),
    1585 => std_logic_vector(to_unsigned(32075, LDPC_TABLE_DATA_WIDTH)),
    1586 => std_logic_vector(to_unsigned(14962, LDPC_TABLE_DATA_WIDTH)),
    1587 => std_logic_vector(to_unsigned(11578, LDPC_TABLE_DATA_WIDTH)),
    1588 => std_logic_vector(to_unsigned(11204, LDPC_TABLE_DATA_WIDTH)),
    1589 => std_logic_vector(to_unsigned(9217, LDPC_TABLE_DATA_WIDTH)),
    1590 => std_logic_vector(to_unsigned(10485, LDPC_TABLE_DATA_WIDTH)),
    1591 => std_logic_vector(to_unsigned(23062, LDPC_TABLE_DATA_WIDTH)),
    1592 => std_logic_vector(to_unsigned(30936, LDPC_TABLE_DATA_WIDTH)),
    1593 => std_logic_vector(to_unsigned(17892, LDPC_TABLE_DATA_WIDTH)),
    1594 => std_logic_vector(to_unsigned(24204, LDPC_TABLE_DATA_WIDTH)),
    1595 => std_logic_vector(to_unsigned(24885, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1596 => std_logic_vector(to_unsigned(32490, LDPC_TABLE_DATA_WIDTH)),
    1597 => std_logic_vector(to_unsigned(18086, LDPC_TABLE_DATA_WIDTH)),
    1598 => std_logic_vector(to_unsigned(18007, LDPC_TABLE_DATA_WIDTH)),
    1599 => std_logic_vector(to_unsigned(4957, LDPC_TABLE_DATA_WIDTH)),
    1600 => std_logic_vector(to_unsigned(7285, LDPC_TABLE_DATA_WIDTH)),
    1601 => std_logic_vector(to_unsigned(32073, LDPC_TABLE_DATA_WIDTH)),
    1602 => std_logic_vector(to_unsigned(19038, LDPC_TABLE_DATA_WIDTH)),
    1603 => std_logic_vector(to_unsigned(7152, LDPC_TABLE_DATA_WIDTH)),
    1604 => std_logic_vector(to_unsigned(12486, LDPC_TABLE_DATA_WIDTH)),
    1605 => std_logic_vector(to_unsigned(13483, LDPC_TABLE_DATA_WIDTH)),
    1606 => std_logic_vector(to_unsigned(24808, LDPC_TABLE_DATA_WIDTH)),
    1607 => std_logic_vector(to_unsigned(21759, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1608 => std_logic_vector(to_unsigned(32321, LDPC_TABLE_DATA_WIDTH)),
    1609 => std_logic_vector(to_unsigned(10839, LDPC_TABLE_DATA_WIDTH)),
    1610 => std_logic_vector(to_unsigned(15620, LDPC_TABLE_DATA_WIDTH)),
    1611 => std_logic_vector(to_unsigned(33521, LDPC_TABLE_DATA_WIDTH)),
    1612 => std_logic_vector(to_unsigned(23030, LDPC_TABLE_DATA_WIDTH)),
    1613 => std_logic_vector(to_unsigned(10646, LDPC_TABLE_DATA_WIDTH)),
    1614 => std_logic_vector(to_unsigned(26236, LDPC_TABLE_DATA_WIDTH)),
    1615 => std_logic_vector(to_unsigned(19744, LDPC_TABLE_DATA_WIDTH)),
    1616 => std_logic_vector(to_unsigned(21713, LDPC_TABLE_DATA_WIDTH)),
    1617 => std_logic_vector(to_unsigned(36784, LDPC_TABLE_DATA_WIDTH)),
    1618 => std_logic_vector(to_unsigned(8016, LDPC_TABLE_DATA_WIDTH)),
    1619 => std_logic_vector(to_unsigned(12869, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1620 => std_logic_vector(to_unsigned(35597, LDPC_TABLE_DATA_WIDTH)),
    1621 => std_logic_vector(to_unsigned(11129, LDPC_TABLE_DATA_WIDTH)),
    1622 => std_logic_vector(to_unsigned(17948, LDPC_TABLE_DATA_WIDTH)),
    1623 => std_logic_vector(to_unsigned(26160, LDPC_TABLE_DATA_WIDTH)),
    1624 => std_logic_vector(to_unsigned(14729, LDPC_TABLE_DATA_WIDTH)),
    1625 => std_logic_vector(to_unsigned(31943, LDPC_TABLE_DATA_WIDTH)),
    1626 => std_logic_vector(to_unsigned(20416, LDPC_TABLE_DATA_WIDTH)),
    1627 => std_logic_vector(to_unsigned(10000, LDPC_TABLE_DATA_WIDTH)),
    1628 => std_logic_vector(to_unsigned(7882, LDPC_TABLE_DATA_WIDTH)),
    1629 => std_logic_vector(to_unsigned(31380, LDPC_TABLE_DATA_WIDTH)),
    1630 => std_logic_vector(to_unsigned(27858, LDPC_TABLE_DATA_WIDTH)),
    1631 => std_logic_vector(to_unsigned(33356, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1632 => std_logic_vector(to_unsigned(14125, LDPC_TABLE_DATA_WIDTH)),
    1633 => std_logic_vector(to_unsigned(12131, LDPC_TABLE_DATA_WIDTH)),
    1634 => std_logic_vector(to_unsigned(36199, LDPC_TABLE_DATA_WIDTH)),
    1635 => std_logic_vector(to_unsigned(4058, LDPC_TABLE_DATA_WIDTH)),
    1636 => std_logic_vector(to_unsigned(35992, LDPC_TABLE_DATA_WIDTH)),
    1637 => std_logic_vector(to_unsigned(36594, LDPC_TABLE_DATA_WIDTH)),
    1638 => std_logic_vector(to_unsigned(33698, LDPC_TABLE_DATA_WIDTH)),
    1639 => std_logic_vector(to_unsigned(15475, LDPC_TABLE_DATA_WIDTH)),
    1640 => std_logic_vector(to_unsigned(1566, LDPC_TABLE_DATA_WIDTH)),
    1641 => std_logic_vector(to_unsigned(18498, LDPC_TABLE_DATA_WIDTH)),
    1642 => std_logic_vector(to_unsigned(12725, LDPC_TABLE_DATA_WIDTH)),
    1643 => std_logic_vector(to_unsigned(7067, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1644 => std_logic_vector(to_unsigned(17406, LDPC_TABLE_DATA_WIDTH)),
    1645 => std_logic_vector(to_unsigned(8372, LDPC_TABLE_DATA_WIDTH)),
    1646 => std_logic_vector(to_unsigned(35437, LDPC_TABLE_DATA_WIDTH)),
    1647 => std_logic_vector(to_unsigned(2888, LDPC_TABLE_DATA_WIDTH)),
    1648 => std_logic_vector(to_unsigned(1184, LDPC_TABLE_DATA_WIDTH)),
    1649 => std_logic_vector(to_unsigned(30068, LDPC_TABLE_DATA_WIDTH)),
    1650 => std_logic_vector(to_unsigned(25802, LDPC_TABLE_DATA_WIDTH)),
    1651 => std_logic_vector(to_unsigned(11056, LDPC_TABLE_DATA_WIDTH)),
    1652 => std_logic_vector(to_unsigned(5507, LDPC_TABLE_DATA_WIDTH)),
    1653 => std_logic_vector(to_unsigned(26313, LDPC_TABLE_DATA_WIDTH)),
    1654 => std_logic_vector(to_unsigned(32205, LDPC_TABLE_DATA_WIDTH)),
    1655 => std_logic_vector(to_unsigned(37232, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1656 => std_logic_vector(to_unsigned(15254, LDPC_TABLE_DATA_WIDTH)),
    1657 => std_logic_vector(to_unsigned(5365, LDPC_TABLE_DATA_WIDTH)),
    1658 => std_logic_vector(to_unsigned(17308, LDPC_TABLE_DATA_WIDTH)),
    1659 => std_logic_vector(to_unsigned(22519, LDPC_TABLE_DATA_WIDTH)),
    1660 => std_logic_vector(to_unsigned(35009, LDPC_TABLE_DATA_WIDTH)),
    1661 => std_logic_vector(to_unsigned(718, LDPC_TABLE_DATA_WIDTH)),
    1662 => std_logic_vector(to_unsigned(5240, LDPC_TABLE_DATA_WIDTH)),
    1663 => std_logic_vector(to_unsigned(16778, LDPC_TABLE_DATA_WIDTH)),
    1664 => std_logic_vector(to_unsigned(23131, LDPC_TABLE_DATA_WIDTH)),
    1665 => std_logic_vector(to_unsigned(24092, LDPC_TABLE_DATA_WIDTH)),
    1666 => std_logic_vector(to_unsigned(20587, LDPC_TABLE_DATA_WIDTH)),
    1667 => std_logic_vector(to_unsigned(33385, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1668 => std_logic_vector(to_unsigned(27455, LDPC_TABLE_DATA_WIDTH)),
    1669 => std_logic_vector(to_unsigned(17602, LDPC_TABLE_DATA_WIDTH)),
    1670 => std_logic_vector(to_unsigned(4590, LDPC_TABLE_DATA_WIDTH)),
    1671 => std_logic_vector(to_unsigned(21767, LDPC_TABLE_DATA_WIDTH)),
    1672 => std_logic_vector(to_unsigned(22266, LDPC_TABLE_DATA_WIDTH)),
    1673 => std_logic_vector(to_unsigned(27357, LDPC_TABLE_DATA_WIDTH)),
    1674 => std_logic_vector(to_unsigned(30400, LDPC_TABLE_DATA_WIDTH)),
    1675 => std_logic_vector(to_unsigned(8732, LDPC_TABLE_DATA_WIDTH)),
    1676 => std_logic_vector(to_unsigned(5596, LDPC_TABLE_DATA_WIDTH)),
    1677 => std_logic_vector(to_unsigned(3060, LDPC_TABLE_DATA_WIDTH)),
    1678 => std_logic_vector(to_unsigned(33703, LDPC_TABLE_DATA_WIDTH)),
    1679 => std_logic_vector(to_unsigned(3596, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1680 => std_logic_vector(to_unsigned(6882, LDPC_TABLE_DATA_WIDTH)),
    1681 => std_logic_vector(to_unsigned(873, LDPC_TABLE_DATA_WIDTH)),
    1682 => std_logic_vector(to_unsigned(10997, LDPC_TABLE_DATA_WIDTH)),
    1683 => std_logic_vector(to_unsigned(24738, LDPC_TABLE_DATA_WIDTH)),
    1684 => std_logic_vector(to_unsigned(20770, LDPC_TABLE_DATA_WIDTH)),
    1685 => std_logic_vector(to_unsigned(10067, LDPC_TABLE_DATA_WIDTH)),
    1686 => std_logic_vector(to_unsigned(13379, LDPC_TABLE_DATA_WIDTH)),
    1687 => std_logic_vector(to_unsigned(27409, LDPC_TABLE_DATA_WIDTH)),
    1688 => std_logic_vector(to_unsigned(25463, LDPC_TABLE_DATA_WIDTH)),
    1689 => std_logic_vector(to_unsigned(2673, LDPC_TABLE_DATA_WIDTH)),
    1690 => std_logic_vector(to_unsigned(6998, LDPC_TABLE_DATA_WIDTH)),
    1691 => std_logic_vector(to_unsigned(31378, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1692 => std_logic_vector(to_unsigned(15181, LDPC_TABLE_DATA_WIDTH)),
    1693 => std_logic_vector(to_unsigned(13645, LDPC_TABLE_DATA_WIDTH)),
    1694 => std_logic_vector(to_unsigned(34501, LDPC_TABLE_DATA_WIDTH)),
    1695 => std_logic_vector(to_unsigned(3393, LDPC_TABLE_DATA_WIDTH)),
    1696 => std_logic_vector(to_unsigned(3840, LDPC_TABLE_DATA_WIDTH)),
    1697 => std_logic_vector(to_unsigned(35227, LDPC_TABLE_DATA_WIDTH)),
    1698 => std_logic_vector(to_unsigned(15562, LDPC_TABLE_DATA_WIDTH)),
    1699 => std_logic_vector(to_unsigned(23615, LDPC_TABLE_DATA_WIDTH)),
    1700 => std_logic_vector(to_unsigned(38342, LDPC_TABLE_DATA_WIDTH)),
    1701 => std_logic_vector(to_unsigned(12139, LDPC_TABLE_DATA_WIDTH)),
    1702 => std_logic_vector(to_unsigned(19471, LDPC_TABLE_DATA_WIDTH)),
    1703 => std_logic_vector(to_unsigned(15483, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1704 => std_logic_vector(to_unsigned(13350, LDPC_TABLE_DATA_WIDTH)),
    1705 => std_logic_vector(to_unsigned(6707, LDPC_TABLE_DATA_WIDTH)),
    1706 => std_logic_vector(to_unsigned(23709, LDPC_TABLE_DATA_WIDTH)),
    1707 => std_logic_vector(to_unsigned(37204, LDPC_TABLE_DATA_WIDTH)),
    1708 => std_logic_vector(to_unsigned(25778, LDPC_TABLE_DATA_WIDTH)),
    1709 => std_logic_vector(to_unsigned(21082, LDPC_TABLE_DATA_WIDTH)),
    1710 => std_logic_vector(to_unsigned(7511, LDPC_TABLE_DATA_WIDTH)),
    1711 => std_logic_vector(to_unsigned(14588, LDPC_TABLE_DATA_WIDTH)),
    1712 => std_logic_vector(to_unsigned(10010, LDPC_TABLE_DATA_WIDTH)),
    1713 => std_logic_vector(to_unsigned(21854, LDPC_TABLE_DATA_WIDTH)),
    1714 => std_logic_vector(to_unsigned(28375, LDPC_TABLE_DATA_WIDTH)),
    1715 => std_logic_vector(to_unsigned(33591, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1716 => std_logic_vector(to_unsigned(12514, LDPC_TABLE_DATA_WIDTH)),
    1717 => std_logic_vector(to_unsigned(4695, LDPC_TABLE_DATA_WIDTH)),
    1718 => std_logic_vector(to_unsigned(37190, LDPC_TABLE_DATA_WIDTH)),
    1719 => std_logic_vector(to_unsigned(21379, LDPC_TABLE_DATA_WIDTH)),
    1720 => std_logic_vector(to_unsigned(18723, LDPC_TABLE_DATA_WIDTH)),
    1721 => std_logic_vector(to_unsigned(5802, LDPC_TABLE_DATA_WIDTH)),
    1722 => std_logic_vector(to_unsigned(7182, LDPC_TABLE_DATA_WIDTH)),
    1723 => std_logic_vector(to_unsigned(2529, LDPC_TABLE_DATA_WIDTH)),
    1724 => std_logic_vector(to_unsigned(29936, LDPC_TABLE_DATA_WIDTH)),
    1725 => std_logic_vector(to_unsigned(35860, LDPC_TABLE_DATA_WIDTH)),
    1726 => std_logic_vector(to_unsigned(28338, LDPC_TABLE_DATA_WIDTH)),
    1727 => std_logic_vector(to_unsigned(10835, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1728 => std_logic_vector(to_unsigned(34283, LDPC_TABLE_DATA_WIDTH)),
    1729 => std_logic_vector(to_unsigned(25610, LDPC_TABLE_DATA_WIDTH)),
    1730 => std_logic_vector(to_unsigned(33026, LDPC_TABLE_DATA_WIDTH)),
    1731 => std_logic_vector(to_unsigned(31017, LDPC_TABLE_DATA_WIDTH)),
    1732 => std_logic_vector(to_unsigned(21259, LDPC_TABLE_DATA_WIDTH)),
    1733 => std_logic_vector(to_unsigned(2165, LDPC_TABLE_DATA_WIDTH)),
    1734 => std_logic_vector(to_unsigned(21807, LDPC_TABLE_DATA_WIDTH)),
    1735 => std_logic_vector(to_unsigned(37578, LDPC_TABLE_DATA_WIDTH)),
    1736 => std_logic_vector(to_unsigned(1175, LDPC_TABLE_DATA_WIDTH)),
    1737 => std_logic_vector(to_unsigned(16710, LDPC_TABLE_DATA_WIDTH)),
    1738 => std_logic_vector(to_unsigned(21939, LDPC_TABLE_DATA_WIDTH)),
    1739 => std_logic_vector(to_unsigned(30841, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1740 => std_logic_vector(to_unsigned(27292, LDPC_TABLE_DATA_WIDTH)),
    1741 => std_logic_vector(to_unsigned(33730, LDPC_TABLE_DATA_WIDTH)),
    1742 => std_logic_vector(to_unsigned(6836, LDPC_TABLE_DATA_WIDTH)),
    1743 => std_logic_vector(to_unsigned(26476, LDPC_TABLE_DATA_WIDTH)),
    1744 => std_logic_vector(to_unsigned(27539, LDPC_TABLE_DATA_WIDTH)),
    1745 => std_logic_vector(to_unsigned(35784, LDPC_TABLE_DATA_WIDTH)),
    1746 => std_logic_vector(to_unsigned(18245, LDPC_TABLE_DATA_WIDTH)),
    1747 => std_logic_vector(to_unsigned(16394, LDPC_TABLE_DATA_WIDTH)),
    1748 => std_logic_vector(to_unsigned(17939, LDPC_TABLE_DATA_WIDTH)),
    1749 => std_logic_vector(to_unsigned(23094, LDPC_TABLE_DATA_WIDTH)),
    1750 => std_logic_vector(to_unsigned(19216, LDPC_TABLE_DATA_WIDTH)),
    1751 => std_logic_vector(to_unsigned(17432, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1752 => std_logic_vector(to_unsigned(11655, LDPC_TABLE_DATA_WIDTH)),
    1753 => std_logic_vector(to_unsigned(6183, LDPC_TABLE_DATA_WIDTH)),
    1754 => std_logic_vector(to_unsigned(38708, LDPC_TABLE_DATA_WIDTH)),
    1755 => std_logic_vector(to_unsigned(28408, LDPC_TABLE_DATA_WIDTH)),
    1756 => std_logic_vector(to_unsigned(35157, LDPC_TABLE_DATA_WIDTH)),
    1757 => std_logic_vector(to_unsigned(17089, LDPC_TABLE_DATA_WIDTH)),
    1758 => std_logic_vector(to_unsigned(13998, LDPC_TABLE_DATA_WIDTH)),
    1759 => std_logic_vector(to_unsigned(36029, LDPC_TABLE_DATA_WIDTH)),
    1760 => std_logic_vector(to_unsigned(15052, LDPC_TABLE_DATA_WIDTH)),
    1761 => std_logic_vector(to_unsigned(16617, LDPC_TABLE_DATA_WIDTH)),
    1762 => std_logic_vector(to_unsigned(5638, LDPC_TABLE_DATA_WIDTH)),
    1763 => std_logic_vector(to_unsigned(36464, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1764 => std_logic_vector(to_unsigned(15693, LDPC_TABLE_DATA_WIDTH)),
    1765 => std_logic_vector(to_unsigned(28923, LDPC_TABLE_DATA_WIDTH)),
    1766 => std_logic_vector(to_unsigned(26245, LDPC_TABLE_DATA_WIDTH)),
    1767 => std_logic_vector(to_unsigned(9432, LDPC_TABLE_DATA_WIDTH)),
    1768 => std_logic_vector(to_unsigned(11675, LDPC_TABLE_DATA_WIDTH)),
    1769 => std_logic_vector(to_unsigned(25720, LDPC_TABLE_DATA_WIDTH)),
    1770 => std_logic_vector(to_unsigned(26405, LDPC_TABLE_DATA_WIDTH)),
    1771 => std_logic_vector(to_unsigned(5838, LDPC_TABLE_DATA_WIDTH)),
    1772 => std_logic_vector(to_unsigned(31851, LDPC_TABLE_DATA_WIDTH)),
    1773 => std_logic_vector(to_unsigned(26898, LDPC_TABLE_DATA_WIDTH)),
    1774 => std_logic_vector(to_unsigned(8090, LDPC_TABLE_DATA_WIDTH)),
    1775 => std_logic_vector(to_unsigned(37037, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1776 => std_logic_vector(to_unsigned(24418, LDPC_TABLE_DATA_WIDTH)),
    1777 => std_logic_vector(to_unsigned(27583, LDPC_TABLE_DATA_WIDTH)),
    1778 => std_logic_vector(to_unsigned(7959, LDPC_TABLE_DATA_WIDTH)),
    1779 => std_logic_vector(to_unsigned(35562, LDPC_TABLE_DATA_WIDTH)),
    1780 => std_logic_vector(to_unsigned(37771, LDPC_TABLE_DATA_WIDTH)),
    1781 => std_logic_vector(to_unsigned(17784, LDPC_TABLE_DATA_WIDTH)),
    1782 => std_logic_vector(to_unsigned(11382, LDPC_TABLE_DATA_WIDTH)),
    1783 => std_logic_vector(to_unsigned(11156, LDPC_TABLE_DATA_WIDTH)),
    1784 => std_logic_vector(to_unsigned(37855, LDPC_TABLE_DATA_WIDTH)),
    1785 => std_logic_vector(to_unsigned(7073, LDPC_TABLE_DATA_WIDTH)),
    1786 => std_logic_vector(to_unsigned(21685, LDPC_TABLE_DATA_WIDTH)),
    1787 => std_logic_vector(to_unsigned(34515, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1788 => std_logic_vector(to_unsigned(10977, LDPC_TABLE_DATA_WIDTH)),
    1789 => std_logic_vector(to_unsigned(13633, LDPC_TABLE_DATA_WIDTH)),
    1790 => std_logic_vector(to_unsigned(30969, LDPC_TABLE_DATA_WIDTH)),
    1791 => std_logic_vector(to_unsigned(7516, LDPC_TABLE_DATA_WIDTH)),
    1792 => std_logic_vector(to_unsigned(11943, LDPC_TABLE_DATA_WIDTH)),
    1793 => std_logic_vector(to_unsigned(18199, LDPC_TABLE_DATA_WIDTH)),
    1794 => std_logic_vector(to_unsigned(5231, LDPC_TABLE_DATA_WIDTH)),
    1795 => std_logic_vector(to_unsigned(13825, LDPC_TABLE_DATA_WIDTH)),
    1796 => std_logic_vector(to_unsigned(19589, LDPC_TABLE_DATA_WIDTH)),
    1797 => std_logic_vector(to_unsigned(23661, LDPC_TABLE_DATA_WIDTH)),
    1798 => std_logic_vector(to_unsigned(11150, LDPC_TABLE_DATA_WIDTH)),
    1799 => std_logic_vector(to_unsigned(35602, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1800 => std_logic_vector(to_unsigned(19124, LDPC_TABLE_DATA_WIDTH)),
    1801 => std_logic_vector(to_unsigned(30774, LDPC_TABLE_DATA_WIDTH)),
    1802 => std_logic_vector(to_unsigned(6670, LDPC_TABLE_DATA_WIDTH)),
    1803 => std_logic_vector(to_unsigned(37344, LDPC_TABLE_DATA_WIDTH)),
    1804 => std_logic_vector(to_unsigned(16510, LDPC_TABLE_DATA_WIDTH)),
    1805 => std_logic_vector(to_unsigned(26317, LDPC_TABLE_DATA_WIDTH)),
    1806 => std_logic_vector(to_unsigned(23518, LDPC_TABLE_DATA_WIDTH)),
    1807 => std_logic_vector(to_unsigned(22957, LDPC_TABLE_DATA_WIDTH)),
    1808 => std_logic_vector(to_unsigned(6348, LDPC_TABLE_DATA_WIDTH)),
    1809 => std_logic_vector(to_unsigned(34069, LDPC_TABLE_DATA_WIDTH)),
    1810 => std_logic_vector(to_unsigned(8845, LDPC_TABLE_DATA_WIDTH)),
    1811 => std_logic_vector(to_unsigned(20175, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1812 => std_logic_vector(to_unsigned(34985, LDPC_TABLE_DATA_WIDTH)),
    1813 => std_logic_vector(to_unsigned(14441, LDPC_TABLE_DATA_WIDTH)),
    1814 => std_logic_vector(to_unsigned(25668, LDPC_TABLE_DATA_WIDTH)),
    1815 => std_logic_vector(to_unsigned(4116, LDPC_TABLE_DATA_WIDTH)),
    1816 => std_logic_vector(to_unsigned(3019, LDPC_TABLE_DATA_WIDTH)),
    1817 => std_logic_vector(to_unsigned(21049, LDPC_TABLE_DATA_WIDTH)),
    1818 => std_logic_vector(to_unsigned(37308, LDPC_TABLE_DATA_WIDTH)),
    1819 => std_logic_vector(to_unsigned(24551, LDPC_TABLE_DATA_WIDTH)),
    1820 => std_logic_vector(to_unsigned(24727, LDPC_TABLE_DATA_WIDTH)),
    1821 => std_logic_vector(to_unsigned(20104, LDPC_TABLE_DATA_WIDTH)),
    1822 => std_logic_vector(to_unsigned(24850, LDPC_TABLE_DATA_WIDTH)),
    1823 => std_logic_vector(to_unsigned(12114, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1824 => std_logic_vector(to_unsigned(38187, LDPC_TABLE_DATA_WIDTH)),
    1825 => std_logic_vector(to_unsigned(28527, LDPC_TABLE_DATA_WIDTH)),
    1826 => std_logic_vector(to_unsigned(13108, LDPC_TABLE_DATA_WIDTH)),
    1827 => std_logic_vector(to_unsigned(13985, LDPC_TABLE_DATA_WIDTH)),
    1828 => std_logic_vector(to_unsigned(1425, LDPC_TABLE_DATA_WIDTH)),
    1829 => std_logic_vector(to_unsigned(21477, LDPC_TABLE_DATA_WIDTH)),
    1830 => std_logic_vector(to_unsigned(30807, LDPC_TABLE_DATA_WIDTH)),
    1831 => std_logic_vector(to_unsigned(8613, LDPC_TABLE_DATA_WIDTH)),
    1832 => std_logic_vector(to_unsigned(26241, LDPC_TABLE_DATA_WIDTH)),
    1833 => std_logic_vector(to_unsigned(33368, LDPC_TABLE_DATA_WIDTH)),
    1834 => std_logic_vector(to_unsigned(35913, LDPC_TABLE_DATA_WIDTH)),
    1835 => std_logic_vector(to_unsigned(32477, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1836 => std_logic_vector(to_unsigned(5903, LDPC_TABLE_DATA_WIDTH)),
    1837 => std_logic_vector(to_unsigned(34390, LDPC_TABLE_DATA_WIDTH)),
    1838 => std_logic_vector(to_unsigned(24641, LDPC_TABLE_DATA_WIDTH)),
    1839 => std_logic_vector(to_unsigned(26556, LDPC_TABLE_DATA_WIDTH)),
    1840 => std_logic_vector(to_unsigned(23007, LDPC_TABLE_DATA_WIDTH)),
    1841 => std_logic_vector(to_unsigned(27305, LDPC_TABLE_DATA_WIDTH)),
    1842 => std_logic_vector(to_unsigned(38247, LDPC_TABLE_DATA_WIDTH)),
    1843 => std_logic_vector(to_unsigned(2621, LDPC_TABLE_DATA_WIDTH)),
    1844 => std_logic_vector(to_unsigned(9122, LDPC_TABLE_DATA_WIDTH)),
    1845 => std_logic_vector(to_unsigned(32806, LDPC_TABLE_DATA_WIDTH)),
    1846 => std_logic_vector(to_unsigned(21554, LDPC_TABLE_DATA_WIDTH)),
    1847 => std_logic_vector(to_unsigned(18685, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1848 => std_logic_vector(to_unsigned(17287, LDPC_TABLE_DATA_WIDTH)),
    1849 => std_logic_vector(to_unsigned(27292, LDPC_TABLE_DATA_WIDTH)),
    1850 => std_logic_vector(to_unsigned(19033, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1851 => std_logic_vector(to_unsigned(25796, LDPC_TABLE_DATA_WIDTH)),
    1852 => std_logic_vector(to_unsigned(31795, LDPC_TABLE_DATA_WIDTH)),
    1853 => std_logic_vector(to_unsigned(12152, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1854 => std_logic_vector(to_unsigned(12184, LDPC_TABLE_DATA_WIDTH)),
    1855 => std_logic_vector(to_unsigned(35088, LDPC_TABLE_DATA_WIDTH)),
    1856 => std_logic_vector(to_unsigned(31226, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1857 => std_logic_vector(to_unsigned(38263, LDPC_TABLE_DATA_WIDTH)),
    1858 => std_logic_vector(to_unsigned(33386, LDPC_TABLE_DATA_WIDTH)),
    1859 => std_logic_vector(to_unsigned(24892, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1860 => std_logic_vector(to_unsigned(23114, LDPC_TABLE_DATA_WIDTH)),
    1861 => std_logic_vector(to_unsigned(37995, LDPC_TABLE_DATA_WIDTH)),
    1862 => std_logic_vector(to_unsigned(29796, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1863 => std_logic_vector(to_unsigned(34336, LDPC_TABLE_DATA_WIDTH)),
    1864 => std_logic_vector(to_unsigned(10551, LDPC_TABLE_DATA_WIDTH)),
    1865 => std_logic_vector(to_unsigned(36245, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1866 => std_logic_vector(to_unsigned(35407, LDPC_TABLE_DATA_WIDTH)),
    1867 => std_logic_vector(to_unsigned(175, LDPC_TABLE_DATA_WIDTH)),
    1868 => std_logic_vector(to_unsigned(7203, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1869 => std_logic_vector(to_unsigned(14654, LDPC_TABLE_DATA_WIDTH)),
    1870 => std_logic_vector(to_unsigned(38201, LDPC_TABLE_DATA_WIDTH)),
    1871 => std_logic_vector(to_unsigned(22605, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1872 => std_logic_vector(to_unsigned(28404, LDPC_TABLE_DATA_WIDTH)),
    1873 => std_logic_vector(to_unsigned(6595, LDPC_TABLE_DATA_WIDTH)),
    1874 => std_logic_vector(to_unsigned(1018, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1875 => std_logic_vector(to_unsigned(19932, LDPC_TABLE_DATA_WIDTH)),
    1876 => std_logic_vector(to_unsigned(3524, LDPC_TABLE_DATA_WIDTH)),
    1877 => std_logic_vector(to_unsigned(29305, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1878 => std_logic_vector(to_unsigned(31749, LDPC_TABLE_DATA_WIDTH)),
    1879 => std_logic_vector(to_unsigned(20247, LDPC_TABLE_DATA_WIDTH)),
    1880 => std_logic_vector(to_unsigned(8128, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1881 => std_logic_vector(to_unsigned(18026, LDPC_TABLE_DATA_WIDTH)),
    1882 => std_logic_vector(to_unsigned(36357, LDPC_TABLE_DATA_WIDTH)),
    1883 => std_logic_vector(to_unsigned(26735, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1884 => std_logic_vector(to_unsigned(7543, LDPC_TABLE_DATA_WIDTH)),
    1885 => std_logic_vector(to_unsigned(29767, LDPC_TABLE_DATA_WIDTH)),
    1886 => std_logic_vector(to_unsigned(13588, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1887 => std_logic_vector(to_unsigned(13333, LDPC_TABLE_DATA_WIDTH)),
    1888 => std_logic_vector(to_unsigned(25965, LDPC_TABLE_DATA_WIDTH)),
    1889 => std_logic_vector(to_unsigned(8463, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1890 => std_logic_vector(to_unsigned(14504, LDPC_TABLE_DATA_WIDTH)),
    1891 => std_logic_vector(to_unsigned(36796, LDPC_TABLE_DATA_WIDTH)),
    1892 => std_logic_vector(to_unsigned(19710, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1893 => std_logic_vector(to_unsigned(4528, LDPC_TABLE_DATA_WIDTH)),
    1894 => std_logic_vector(to_unsigned(25299, LDPC_TABLE_DATA_WIDTH)),
    1895 => std_logic_vector(to_unsigned(7318, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1896 => std_logic_vector(to_unsigned(35091, LDPC_TABLE_DATA_WIDTH)),
    1897 => std_logic_vector(to_unsigned(25550, LDPC_TABLE_DATA_WIDTH)),
    1898 => std_logic_vector(to_unsigned(14798, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1899 => std_logic_vector(to_unsigned(7824, LDPC_TABLE_DATA_WIDTH)),
    1900 => std_logic_vector(to_unsigned(215, LDPC_TABLE_DATA_WIDTH)),
    1901 => std_logic_vector(to_unsigned(1248, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1902 => std_logic_vector(to_unsigned(30848, LDPC_TABLE_DATA_WIDTH)),
    1903 => std_logic_vector(to_unsigned(5362, LDPC_TABLE_DATA_WIDTH)),
    1904 => std_logic_vector(to_unsigned(17291, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1905 => std_logic_vector(to_unsigned(28932, LDPC_TABLE_DATA_WIDTH)),
    1906 => std_logic_vector(to_unsigned(30249, LDPC_TABLE_DATA_WIDTH)),
    1907 => std_logic_vector(to_unsigned(27073, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1908 => std_logic_vector(to_unsigned(13062, LDPC_TABLE_DATA_WIDTH)),
    1909 => std_logic_vector(to_unsigned(2103, LDPC_TABLE_DATA_WIDTH)),
    1910 => std_logic_vector(to_unsigned(16206, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1911 => std_logic_vector(to_unsigned(7129, LDPC_TABLE_DATA_WIDTH)),
    1912 => std_logic_vector(to_unsigned(32062, LDPC_TABLE_DATA_WIDTH)),
    1913 => std_logic_vector(to_unsigned(19612, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1914 => std_logic_vector(to_unsigned(9512, LDPC_TABLE_DATA_WIDTH)),
    1915 => std_logic_vector(to_unsigned(21936, LDPC_TABLE_DATA_WIDTH)),
    1916 => std_logic_vector(to_unsigned(38833, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1917 => std_logic_vector(to_unsigned(35849, LDPC_TABLE_DATA_WIDTH)),
    1918 => std_logic_vector(to_unsigned(33754, LDPC_TABLE_DATA_WIDTH)),
    1919 => std_logic_vector(to_unsigned(23450, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1920 => std_logic_vector(to_unsigned(18705, LDPC_TABLE_DATA_WIDTH)),
    1921 => std_logic_vector(to_unsigned(28656, LDPC_TABLE_DATA_WIDTH)),
    1922 => std_logic_vector(to_unsigned(18111, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1923 => std_logic_vector(to_unsigned(22749, LDPC_TABLE_DATA_WIDTH)),
    1924 => std_logic_vector(to_unsigned(27456, LDPC_TABLE_DATA_WIDTH)),
    1925 => std_logic_vector(to_unsigned(32187, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1926 => std_logic_vector(to_unsigned(28229, LDPC_TABLE_DATA_WIDTH)),
    1927 => std_logic_vector(to_unsigned(31684, LDPC_TABLE_DATA_WIDTH)),
    1928 => std_logic_vector(to_unsigned(30160, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1929 => std_logic_vector(to_unsigned(15293, LDPC_TABLE_DATA_WIDTH)),
    1930 => std_logic_vector(to_unsigned(8483, LDPC_TABLE_DATA_WIDTH)),
    1931 => std_logic_vector(to_unsigned(28002, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1932 => std_logic_vector(to_unsigned(14880, LDPC_TABLE_DATA_WIDTH)),
    1933 => std_logic_vector(to_unsigned(13334, LDPC_TABLE_DATA_WIDTH)),
    1934 => std_logic_vector(to_unsigned(12584, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1935 => std_logic_vector(to_unsigned(28646, LDPC_TABLE_DATA_WIDTH)),
    1936 => std_logic_vector(to_unsigned(2558, LDPC_TABLE_DATA_WIDTH)),
    1937 => std_logic_vector(to_unsigned(19687, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1938 => std_logic_vector(to_unsigned(6259, LDPC_TABLE_DATA_WIDTH)),
    1939 => std_logic_vector(to_unsigned(4499, LDPC_TABLE_DATA_WIDTH)),
    1940 => std_logic_vector(to_unsigned(26336, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1941 => std_logic_vector(to_unsigned(11952, LDPC_TABLE_DATA_WIDTH)),
    1942 => std_logic_vector(to_unsigned(28386, LDPC_TABLE_DATA_WIDTH)),
    1943 => std_logic_vector(to_unsigned(8405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1944 => std_logic_vector(to_unsigned(10609, LDPC_TABLE_DATA_WIDTH)),
    1945 => std_logic_vector(to_unsigned(961, LDPC_TABLE_DATA_WIDTH)),
    1946 => std_logic_vector(to_unsigned(7582, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1947 => std_logic_vector(to_unsigned(10423, LDPC_TABLE_DATA_WIDTH)),
    1948 => std_logic_vector(to_unsigned(13191, LDPC_TABLE_DATA_WIDTH)),
    1949 => std_logic_vector(to_unsigned(26818, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1950 => std_logic_vector(to_unsigned(15922, LDPC_TABLE_DATA_WIDTH)),
    1951 => std_logic_vector(to_unsigned(36654, LDPC_TABLE_DATA_WIDTH)),
    1952 => std_logic_vector(to_unsigned(21450, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1953 => std_logic_vector(to_unsigned(10492, LDPC_TABLE_DATA_WIDTH)),
    1954 => std_logic_vector(to_unsigned(1532, LDPC_TABLE_DATA_WIDTH)),
    1955 => std_logic_vector(to_unsigned(1205, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1956 => std_logic_vector(to_unsigned(30551, LDPC_TABLE_DATA_WIDTH)),
    1957 => std_logic_vector(to_unsigned(36482, LDPC_TABLE_DATA_WIDTH)),
    1958 => std_logic_vector(to_unsigned(22153, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1959 => std_logic_vector(to_unsigned(5156, LDPC_TABLE_DATA_WIDTH)),
    1960 => std_logic_vector(to_unsigned(11330, LDPC_TABLE_DATA_WIDTH)),
    1961 => std_logic_vector(to_unsigned(34243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1962 => std_logic_vector(to_unsigned(28616, LDPC_TABLE_DATA_WIDTH)),
    1963 => std_logic_vector(to_unsigned(35369, LDPC_TABLE_DATA_WIDTH)),
    1964 => std_logic_vector(to_unsigned(13322, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1965 => std_logic_vector(to_unsigned(8962, LDPC_TABLE_DATA_WIDTH)),
    1966 => std_logic_vector(to_unsigned(1485, LDPC_TABLE_DATA_WIDTH)),
    1967 => std_logic_vector(to_unsigned(21186, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1968 => std_logic_vector(to_unsigned(23541, LDPC_TABLE_DATA_WIDTH)),
    1969 => std_logic_vector(to_unsigned(17445, LDPC_TABLE_DATA_WIDTH)),
    1970 => std_logic_vector(to_unsigned(35561, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1971 => std_logic_vector(to_unsigned(33133, LDPC_TABLE_DATA_WIDTH)),
    1972 => std_logic_vector(to_unsigned(11593, LDPC_TABLE_DATA_WIDTH)),
    1973 => std_logic_vector(to_unsigned(19895, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1974 => std_logic_vector(to_unsigned(33917, LDPC_TABLE_DATA_WIDTH)),
    1975 => std_logic_vector(to_unsigned(7863, LDPC_TABLE_DATA_WIDTH)),
    1976 => std_logic_vector(to_unsigned(33651, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1977 => std_logic_vector(to_unsigned(20063, LDPC_TABLE_DATA_WIDTH)),
    1978 => std_logic_vector(to_unsigned(28331, LDPC_TABLE_DATA_WIDTH)),
    1979 => std_logic_vector(to_unsigned(10702, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1980 => std_logic_vector(to_unsigned(13195, LDPC_TABLE_DATA_WIDTH)),
    1981 => std_logic_vector(to_unsigned(21107, LDPC_TABLE_DATA_WIDTH)),
    1982 => std_logic_vector(to_unsigned(21859, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1983 => std_logic_vector(to_unsigned(4364, LDPC_TABLE_DATA_WIDTH)),
    1984 => std_logic_vector(to_unsigned(31137, LDPC_TABLE_DATA_WIDTH)),
    1985 => std_logic_vector(to_unsigned(4804, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1986 => std_logic_vector(to_unsigned(5585, LDPC_TABLE_DATA_WIDTH)),
    1987 => std_logic_vector(to_unsigned(2037, LDPC_TABLE_DATA_WIDTH)),
    1988 => std_logic_vector(to_unsigned(4830, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    1989 => std_logic_vector(to_unsigned(30672, LDPC_TABLE_DATA_WIDTH)),
    1990 => std_logic_vector(to_unsigned(16927, LDPC_TABLE_DATA_WIDTH)),
    1991 => std_logic_vector(to_unsigned(14800, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C3_4
    1992 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    1993 => std_logic_vector(to_unsigned(6385, LDPC_TABLE_DATA_WIDTH)),
    1994 => std_logic_vector(to_unsigned(7901, LDPC_TABLE_DATA_WIDTH)),
    1995 => std_logic_vector(to_unsigned(14611, LDPC_TABLE_DATA_WIDTH)),
    1996 => std_logic_vector(to_unsigned(13389, LDPC_TABLE_DATA_WIDTH)),
    1997 => std_logic_vector(to_unsigned(11200, LDPC_TABLE_DATA_WIDTH)),
    1998 => std_logic_vector(to_unsigned(3252, LDPC_TABLE_DATA_WIDTH)),
    1999 => std_logic_vector(to_unsigned(5243, LDPC_TABLE_DATA_WIDTH)),
    2000 => std_logic_vector(to_unsigned(2504, LDPC_TABLE_DATA_WIDTH)),
    2001 => std_logic_vector(to_unsigned(2722, LDPC_TABLE_DATA_WIDTH)),
    2002 => std_logic_vector(to_unsigned(821, LDPC_TABLE_DATA_WIDTH)),
    2003 => std_logic_vector(to_unsigned(7374, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2004 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    2005 => std_logic_vector(to_unsigned(11359, LDPC_TABLE_DATA_WIDTH)),
    2006 => std_logic_vector(to_unsigned(2698, LDPC_TABLE_DATA_WIDTH)),
    2007 => std_logic_vector(to_unsigned(357, LDPC_TABLE_DATA_WIDTH)),
    2008 => std_logic_vector(to_unsigned(13824, LDPC_TABLE_DATA_WIDTH)),
    2009 => std_logic_vector(to_unsigned(12772, LDPC_TABLE_DATA_WIDTH)),
    2010 => std_logic_vector(to_unsigned(7244, LDPC_TABLE_DATA_WIDTH)),
    2011 => std_logic_vector(to_unsigned(6752, LDPC_TABLE_DATA_WIDTH)),
    2012 => std_logic_vector(to_unsigned(15310, LDPC_TABLE_DATA_WIDTH)),
    2013 => std_logic_vector(to_unsigned(852, LDPC_TABLE_DATA_WIDTH)),
    2014 => std_logic_vector(to_unsigned(2001, LDPC_TABLE_DATA_WIDTH)),
    2015 => std_logic_vector(to_unsigned(11417, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2016 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    2017 => std_logic_vector(to_unsigned(7862, LDPC_TABLE_DATA_WIDTH)),
    2018 => std_logic_vector(to_unsigned(7977, LDPC_TABLE_DATA_WIDTH)),
    2019 => std_logic_vector(to_unsigned(6321, LDPC_TABLE_DATA_WIDTH)),
    2020 => std_logic_vector(to_unsigned(13612, LDPC_TABLE_DATA_WIDTH)),
    2021 => std_logic_vector(to_unsigned(12197, LDPC_TABLE_DATA_WIDTH)),
    2022 => std_logic_vector(to_unsigned(14449, LDPC_TABLE_DATA_WIDTH)),
    2023 => std_logic_vector(to_unsigned(15137, LDPC_TABLE_DATA_WIDTH)),
    2024 => std_logic_vector(to_unsigned(13860, LDPC_TABLE_DATA_WIDTH)),
    2025 => std_logic_vector(to_unsigned(1708, LDPC_TABLE_DATA_WIDTH)),
    2026 => std_logic_vector(to_unsigned(6399, LDPC_TABLE_DATA_WIDTH)),
    2027 => std_logic_vector(to_unsigned(13444, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2028 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    2029 => std_logic_vector(to_unsigned(1560, LDPC_TABLE_DATA_WIDTH)),
    2030 => std_logic_vector(to_unsigned(11804, LDPC_TABLE_DATA_WIDTH)),
    2031 => std_logic_vector(to_unsigned(6975, LDPC_TABLE_DATA_WIDTH)),
    2032 => std_logic_vector(to_unsigned(13292, LDPC_TABLE_DATA_WIDTH)),
    2033 => std_logic_vector(to_unsigned(3646, LDPC_TABLE_DATA_WIDTH)),
    2034 => std_logic_vector(to_unsigned(3812, LDPC_TABLE_DATA_WIDTH)),
    2035 => std_logic_vector(to_unsigned(8772, LDPC_TABLE_DATA_WIDTH)),
    2036 => std_logic_vector(to_unsigned(7306, LDPC_TABLE_DATA_WIDTH)),
    2037 => std_logic_vector(to_unsigned(5795, LDPC_TABLE_DATA_WIDTH)),
    2038 => std_logic_vector(to_unsigned(14327, LDPC_TABLE_DATA_WIDTH)),
    2039 => std_logic_vector(to_unsigned(7866, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2040 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    2041 => std_logic_vector(to_unsigned(7626, LDPC_TABLE_DATA_WIDTH)),
    2042 => std_logic_vector(to_unsigned(11407, LDPC_TABLE_DATA_WIDTH)),
    2043 => std_logic_vector(to_unsigned(14599, LDPC_TABLE_DATA_WIDTH)),
    2044 => std_logic_vector(to_unsigned(9689, LDPC_TABLE_DATA_WIDTH)),
    2045 => std_logic_vector(to_unsigned(1628, LDPC_TABLE_DATA_WIDTH)),
    2046 => std_logic_vector(to_unsigned(2113, LDPC_TABLE_DATA_WIDTH)),
    2047 => std_logic_vector(to_unsigned(10809, LDPC_TABLE_DATA_WIDTH)),
    2048 => std_logic_vector(to_unsigned(9283, LDPC_TABLE_DATA_WIDTH)),
    2049 => std_logic_vector(to_unsigned(1230, LDPC_TABLE_DATA_WIDTH)),
    2050 => std_logic_vector(to_unsigned(15241, LDPC_TABLE_DATA_WIDTH)),
    2051 => std_logic_vector(to_unsigned(4870, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2052 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    2053 => std_logic_vector(to_unsigned(1610, LDPC_TABLE_DATA_WIDTH)),
    2054 => std_logic_vector(to_unsigned(5699, LDPC_TABLE_DATA_WIDTH)),
    2055 => std_logic_vector(to_unsigned(15876, LDPC_TABLE_DATA_WIDTH)),
    2056 => std_logic_vector(to_unsigned(9446, LDPC_TABLE_DATA_WIDTH)),
    2057 => std_logic_vector(to_unsigned(12515, LDPC_TABLE_DATA_WIDTH)),
    2058 => std_logic_vector(to_unsigned(1400, LDPC_TABLE_DATA_WIDTH)),
    2059 => std_logic_vector(to_unsigned(6303, LDPC_TABLE_DATA_WIDTH)),
    2060 => std_logic_vector(to_unsigned(5411, LDPC_TABLE_DATA_WIDTH)),
    2061 => std_logic_vector(to_unsigned(14181, LDPC_TABLE_DATA_WIDTH)),
    2062 => std_logic_vector(to_unsigned(13925, LDPC_TABLE_DATA_WIDTH)),
    2063 => std_logic_vector(to_unsigned(7358, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2064 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    2065 => std_logic_vector(to_unsigned(4059, LDPC_TABLE_DATA_WIDTH)),
    2066 => std_logic_vector(to_unsigned(8836, LDPC_TABLE_DATA_WIDTH)),
    2067 => std_logic_vector(to_unsigned(3405, LDPC_TABLE_DATA_WIDTH)),
    2068 => std_logic_vector(to_unsigned(7853, LDPC_TABLE_DATA_WIDTH)),
    2069 => std_logic_vector(to_unsigned(7992, LDPC_TABLE_DATA_WIDTH)),
    2070 => std_logic_vector(to_unsigned(15336, LDPC_TABLE_DATA_WIDTH)),
    2071 => std_logic_vector(to_unsigned(5970, LDPC_TABLE_DATA_WIDTH)),
    2072 => std_logic_vector(to_unsigned(10368, LDPC_TABLE_DATA_WIDTH)),
    2073 => std_logic_vector(to_unsigned(10278, LDPC_TABLE_DATA_WIDTH)),
    2074 => std_logic_vector(to_unsigned(9675, LDPC_TABLE_DATA_WIDTH)),
    2075 => std_logic_vector(to_unsigned(4651, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2076 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    2077 => std_logic_vector(to_unsigned(4441, LDPC_TABLE_DATA_WIDTH)),
    2078 => std_logic_vector(to_unsigned(3963, LDPC_TABLE_DATA_WIDTH)),
    2079 => std_logic_vector(to_unsigned(9153, LDPC_TABLE_DATA_WIDTH)),
    2080 => std_logic_vector(to_unsigned(2109, LDPC_TABLE_DATA_WIDTH)),
    2081 => std_logic_vector(to_unsigned(12683, LDPC_TABLE_DATA_WIDTH)),
    2082 => std_logic_vector(to_unsigned(7459, LDPC_TABLE_DATA_WIDTH)),
    2083 => std_logic_vector(to_unsigned(12030, LDPC_TABLE_DATA_WIDTH)),
    2084 => std_logic_vector(to_unsigned(12221, LDPC_TABLE_DATA_WIDTH)),
    2085 => std_logic_vector(to_unsigned(629, LDPC_TABLE_DATA_WIDTH)),
    2086 => std_logic_vector(to_unsigned(15212, LDPC_TABLE_DATA_WIDTH)),
    2087 => std_logic_vector(to_unsigned(406, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2088 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    2089 => std_logic_vector(to_unsigned(6007, LDPC_TABLE_DATA_WIDTH)),
    2090 => std_logic_vector(to_unsigned(8411, LDPC_TABLE_DATA_WIDTH)),
    2091 => std_logic_vector(to_unsigned(5771, LDPC_TABLE_DATA_WIDTH)),
    2092 => std_logic_vector(to_unsigned(3497, LDPC_TABLE_DATA_WIDTH)),
    2093 => std_logic_vector(to_unsigned(543, LDPC_TABLE_DATA_WIDTH)),
    2094 => std_logic_vector(to_unsigned(14202, LDPC_TABLE_DATA_WIDTH)),
    2095 => std_logic_vector(to_unsigned(875, LDPC_TABLE_DATA_WIDTH)),
    2096 => std_logic_vector(to_unsigned(9186, LDPC_TABLE_DATA_WIDTH)),
    2097 => std_logic_vector(to_unsigned(6235, LDPC_TABLE_DATA_WIDTH)),
    2098 => std_logic_vector(to_unsigned(13908, LDPC_TABLE_DATA_WIDTH)),
    2099 => std_logic_vector(to_unsigned(3563, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2100 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    2101 => std_logic_vector(to_unsigned(3232, LDPC_TABLE_DATA_WIDTH)),
    2102 => std_logic_vector(to_unsigned(6625, LDPC_TABLE_DATA_WIDTH)),
    2103 => std_logic_vector(to_unsigned(4795, LDPC_TABLE_DATA_WIDTH)),
    2104 => std_logic_vector(to_unsigned(546, LDPC_TABLE_DATA_WIDTH)),
    2105 => std_logic_vector(to_unsigned(9781, LDPC_TABLE_DATA_WIDTH)),
    2106 => std_logic_vector(to_unsigned(2071, LDPC_TABLE_DATA_WIDTH)),
    2107 => std_logic_vector(to_unsigned(7312, LDPC_TABLE_DATA_WIDTH)),
    2108 => std_logic_vector(to_unsigned(3399, LDPC_TABLE_DATA_WIDTH)),
    2109 => std_logic_vector(to_unsigned(7250, LDPC_TABLE_DATA_WIDTH)),
    2110 => std_logic_vector(to_unsigned(4932, LDPC_TABLE_DATA_WIDTH)),
    2111 => std_logic_vector(to_unsigned(12652, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2112 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    2113 => std_logic_vector(to_unsigned(8820, LDPC_TABLE_DATA_WIDTH)),
    2114 => std_logic_vector(to_unsigned(10088, LDPC_TABLE_DATA_WIDTH)),
    2115 => std_logic_vector(to_unsigned(11090, LDPC_TABLE_DATA_WIDTH)),
    2116 => std_logic_vector(to_unsigned(7069, LDPC_TABLE_DATA_WIDTH)),
    2117 => std_logic_vector(to_unsigned(6585, LDPC_TABLE_DATA_WIDTH)),
    2118 => std_logic_vector(to_unsigned(13134, LDPC_TABLE_DATA_WIDTH)),
    2119 => std_logic_vector(to_unsigned(10158, LDPC_TABLE_DATA_WIDTH)),
    2120 => std_logic_vector(to_unsigned(7183, LDPC_TABLE_DATA_WIDTH)),
    2121 => std_logic_vector(to_unsigned(488, LDPC_TABLE_DATA_WIDTH)),
    2122 => std_logic_vector(to_unsigned(7455, LDPC_TABLE_DATA_WIDTH)),
    2123 => std_logic_vector(to_unsigned(9238, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2124 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    2125 => std_logic_vector(to_unsigned(1903, LDPC_TABLE_DATA_WIDTH)),
    2126 => std_logic_vector(to_unsigned(10818, LDPC_TABLE_DATA_WIDTH)),
    2127 => std_logic_vector(to_unsigned(119, LDPC_TABLE_DATA_WIDTH)),
    2128 => std_logic_vector(to_unsigned(215, LDPC_TABLE_DATA_WIDTH)),
    2129 => std_logic_vector(to_unsigned(7558, LDPC_TABLE_DATA_WIDTH)),
    2130 => std_logic_vector(to_unsigned(11046, LDPC_TABLE_DATA_WIDTH)),
    2131 => std_logic_vector(to_unsigned(10615, LDPC_TABLE_DATA_WIDTH)),
    2132 => std_logic_vector(to_unsigned(11545, LDPC_TABLE_DATA_WIDTH)),
    2133 => std_logic_vector(to_unsigned(14784, LDPC_TABLE_DATA_WIDTH)),
    2134 => std_logic_vector(to_unsigned(7961, LDPC_TABLE_DATA_WIDTH)),
    2135 => std_logic_vector(to_unsigned(15619, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2136 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    2137 => std_logic_vector(to_unsigned(3655, LDPC_TABLE_DATA_WIDTH)),
    2138 => std_logic_vector(to_unsigned(8736, LDPC_TABLE_DATA_WIDTH)),
    2139 => std_logic_vector(to_unsigned(4917, LDPC_TABLE_DATA_WIDTH)),
    2140 => std_logic_vector(to_unsigned(15874, LDPC_TABLE_DATA_WIDTH)),
    2141 => std_logic_vector(to_unsigned(5129, LDPC_TABLE_DATA_WIDTH)),
    2142 => std_logic_vector(to_unsigned(2134, LDPC_TABLE_DATA_WIDTH)),
    2143 => std_logic_vector(to_unsigned(15944, LDPC_TABLE_DATA_WIDTH)),
    2144 => std_logic_vector(to_unsigned(14768, LDPC_TABLE_DATA_WIDTH)),
    2145 => std_logic_vector(to_unsigned(7150, LDPC_TABLE_DATA_WIDTH)),
    2146 => std_logic_vector(to_unsigned(2692, LDPC_TABLE_DATA_WIDTH)),
    2147 => std_logic_vector(to_unsigned(1469, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2148 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    2149 => std_logic_vector(to_unsigned(8316, LDPC_TABLE_DATA_WIDTH)),
    2150 => std_logic_vector(to_unsigned(3820, LDPC_TABLE_DATA_WIDTH)),
    2151 => std_logic_vector(to_unsigned(505, LDPC_TABLE_DATA_WIDTH)),
    2152 => std_logic_vector(to_unsigned(8923, LDPC_TABLE_DATA_WIDTH)),
    2153 => std_logic_vector(to_unsigned(6757, LDPC_TABLE_DATA_WIDTH)),
    2154 => std_logic_vector(to_unsigned(806, LDPC_TABLE_DATA_WIDTH)),
    2155 => std_logic_vector(to_unsigned(7957, LDPC_TABLE_DATA_WIDTH)),
    2156 => std_logic_vector(to_unsigned(4216, LDPC_TABLE_DATA_WIDTH)),
    2157 => std_logic_vector(to_unsigned(15589, LDPC_TABLE_DATA_WIDTH)),
    2158 => std_logic_vector(to_unsigned(13244, LDPC_TABLE_DATA_WIDTH)),
    2159 => std_logic_vector(to_unsigned(2622, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2160 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    2161 => std_logic_vector(to_unsigned(14463, LDPC_TABLE_DATA_WIDTH)),
    2162 => std_logic_vector(to_unsigned(4852, LDPC_TABLE_DATA_WIDTH)),
    2163 => std_logic_vector(to_unsigned(15733, LDPC_TABLE_DATA_WIDTH)),
    2164 => std_logic_vector(to_unsigned(3041, LDPC_TABLE_DATA_WIDTH)),
    2165 => std_logic_vector(to_unsigned(11193, LDPC_TABLE_DATA_WIDTH)),
    2166 => std_logic_vector(to_unsigned(12860, LDPC_TABLE_DATA_WIDTH)),
    2167 => std_logic_vector(to_unsigned(13673, LDPC_TABLE_DATA_WIDTH)),
    2168 => std_logic_vector(to_unsigned(8152, LDPC_TABLE_DATA_WIDTH)),
    2169 => std_logic_vector(to_unsigned(6551, LDPC_TABLE_DATA_WIDTH)),
    2170 => std_logic_vector(to_unsigned(15108, LDPC_TABLE_DATA_WIDTH)),
    2171 => std_logic_vector(to_unsigned(8758, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2172 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    2173 => std_logic_vector(to_unsigned(3149, LDPC_TABLE_DATA_WIDTH)),
    2174 => std_logic_vector(to_unsigned(11981, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2175 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    2176 => std_logic_vector(to_unsigned(13416, LDPC_TABLE_DATA_WIDTH)),
    2177 => std_logic_vector(to_unsigned(6906, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2178 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    2179 => std_logic_vector(to_unsigned(13098, LDPC_TABLE_DATA_WIDTH)),
    2180 => std_logic_vector(to_unsigned(13352, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2181 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    2182 => std_logic_vector(to_unsigned(2009, LDPC_TABLE_DATA_WIDTH)),
    2183 => std_logic_vector(to_unsigned(14460, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2184 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    2185 => std_logic_vector(to_unsigned(7207, LDPC_TABLE_DATA_WIDTH)),
    2186 => std_logic_vector(to_unsigned(4314, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2187 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    2188 => std_logic_vector(to_unsigned(3312, LDPC_TABLE_DATA_WIDTH)),
    2189 => std_logic_vector(to_unsigned(3945, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2190 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    2191 => std_logic_vector(to_unsigned(4418, LDPC_TABLE_DATA_WIDTH)),
    2192 => std_logic_vector(to_unsigned(6248, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2193 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    2194 => std_logic_vector(to_unsigned(2669, LDPC_TABLE_DATA_WIDTH)),
    2195 => std_logic_vector(to_unsigned(13975, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2196 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    2197 => std_logic_vector(to_unsigned(7571, LDPC_TABLE_DATA_WIDTH)),
    2198 => std_logic_vector(to_unsigned(9023, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2199 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    2200 => std_logic_vector(to_unsigned(14172, LDPC_TABLE_DATA_WIDTH)),
    2201 => std_logic_vector(to_unsigned(2967, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2202 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    2203 => std_logic_vector(to_unsigned(7271, LDPC_TABLE_DATA_WIDTH)),
    2204 => std_logic_vector(to_unsigned(7138, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2205 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    2206 => std_logic_vector(to_unsigned(6135, LDPC_TABLE_DATA_WIDTH)),
    2207 => std_logic_vector(to_unsigned(13670, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2208 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    2209 => std_logic_vector(to_unsigned(7490, LDPC_TABLE_DATA_WIDTH)),
    2210 => std_logic_vector(to_unsigned(14559, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2211 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    2212 => std_logic_vector(to_unsigned(8657, LDPC_TABLE_DATA_WIDTH)),
    2213 => std_logic_vector(to_unsigned(2466, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2214 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    2215 => std_logic_vector(to_unsigned(8599, LDPC_TABLE_DATA_WIDTH)),
    2216 => std_logic_vector(to_unsigned(12834, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2217 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    2218 => std_logic_vector(to_unsigned(3470, LDPC_TABLE_DATA_WIDTH)),
    2219 => std_logic_vector(to_unsigned(3152, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2220 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    2221 => std_logic_vector(to_unsigned(13917, LDPC_TABLE_DATA_WIDTH)),
    2222 => std_logic_vector(to_unsigned(4365, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2223 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    2224 => std_logic_vector(to_unsigned(6024, LDPC_TABLE_DATA_WIDTH)),
    2225 => std_logic_vector(to_unsigned(13730, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2226 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    2227 => std_logic_vector(to_unsigned(10973, LDPC_TABLE_DATA_WIDTH)),
    2228 => std_logic_vector(to_unsigned(14182, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2229 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    2230 => std_logic_vector(to_unsigned(2464, LDPC_TABLE_DATA_WIDTH)),
    2231 => std_logic_vector(to_unsigned(13167, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2232 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    2233 => std_logic_vector(to_unsigned(5281, LDPC_TABLE_DATA_WIDTH)),
    2234 => std_logic_vector(to_unsigned(15049, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2235 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    2236 => std_logic_vector(to_unsigned(1103, LDPC_TABLE_DATA_WIDTH)),
    2237 => std_logic_vector(to_unsigned(1849, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2238 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    2239 => std_logic_vector(to_unsigned(2058, LDPC_TABLE_DATA_WIDTH)),
    2240 => std_logic_vector(to_unsigned(1069, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2241 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    2242 => std_logic_vector(to_unsigned(9654, LDPC_TABLE_DATA_WIDTH)),
    2243 => std_logic_vector(to_unsigned(6095, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2244 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    2245 => std_logic_vector(to_unsigned(14311, LDPC_TABLE_DATA_WIDTH)),
    2246 => std_logic_vector(to_unsigned(7667, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2247 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    2248 => std_logic_vector(to_unsigned(15617, LDPC_TABLE_DATA_WIDTH)),
    2249 => std_logic_vector(to_unsigned(8146, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2250 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    2251 => std_logic_vector(to_unsigned(4588, LDPC_TABLE_DATA_WIDTH)),
    2252 => std_logic_vector(to_unsigned(11218, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2253 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    2254 => std_logic_vector(to_unsigned(13660, LDPC_TABLE_DATA_WIDTH)),
    2255 => std_logic_vector(to_unsigned(6243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2256 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    2257 => std_logic_vector(to_unsigned(8578, LDPC_TABLE_DATA_WIDTH)),
    2258 => std_logic_vector(to_unsigned(7874, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2259 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    2260 => std_logic_vector(to_unsigned(11741, LDPC_TABLE_DATA_WIDTH)),
    2261 => std_logic_vector(to_unsigned(2686, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2262 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    2263 => std_logic_vector(to_unsigned(1022, LDPC_TABLE_DATA_WIDTH)),
    2264 => std_logic_vector(to_unsigned(1264, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2265 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    2266 => std_logic_vector(to_unsigned(12604, LDPC_TABLE_DATA_WIDTH)),
    2267 => std_logic_vector(to_unsigned(9965, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2268 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    2269 => std_logic_vector(to_unsigned(8217, LDPC_TABLE_DATA_WIDTH)),
    2270 => std_logic_vector(to_unsigned(2707, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2271 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    2272 => std_logic_vector(to_unsigned(3156, LDPC_TABLE_DATA_WIDTH)),
    2273 => std_logic_vector(to_unsigned(11793, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2274 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    2275 => std_logic_vector(to_unsigned(354, LDPC_TABLE_DATA_WIDTH)),
    2276 => std_logic_vector(to_unsigned(1514, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2277 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    2278 => std_logic_vector(to_unsigned(6978, LDPC_TABLE_DATA_WIDTH)),
    2279 => std_logic_vector(to_unsigned(14058, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2280 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    2281 => std_logic_vector(to_unsigned(7922, LDPC_TABLE_DATA_WIDTH)),
    2282 => std_logic_vector(to_unsigned(16079, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2283 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    2284 => std_logic_vector(to_unsigned(15087, LDPC_TABLE_DATA_WIDTH)),
    2285 => std_logic_vector(to_unsigned(12138, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2286 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    2287 => std_logic_vector(to_unsigned(5053, LDPC_TABLE_DATA_WIDTH)),
    2288 => std_logic_vector(to_unsigned(6470, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2289 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    2290 => std_logic_vector(to_unsigned(12687, LDPC_TABLE_DATA_WIDTH)),
    2291 => std_logic_vector(to_unsigned(14932, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2292 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    2293 => std_logic_vector(to_unsigned(15458, LDPC_TABLE_DATA_WIDTH)),
    2294 => std_logic_vector(to_unsigned(1763, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2295 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    2296 => std_logic_vector(to_unsigned(8121, LDPC_TABLE_DATA_WIDTH)),
    2297 => std_logic_vector(to_unsigned(1721, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2298 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    2299 => std_logic_vector(to_unsigned(12431, LDPC_TABLE_DATA_WIDTH)),
    2300 => std_logic_vector(to_unsigned(549, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2301 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    2302 => std_logic_vector(to_unsigned(4129, LDPC_TABLE_DATA_WIDTH)),
    2303 => std_logic_vector(to_unsigned(7091, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2304 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    2305 => std_logic_vector(to_unsigned(1426, LDPC_TABLE_DATA_WIDTH)),
    2306 => std_logic_vector(to_unsigned(8415, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2307 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    2308 => std_logic_vector(to_unsigned(9783, LDPC_TABLE_DATA_WIDTH)),
    2309 => std_logic_vector(to_unsigned(7604, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2310 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    2311 => std_logic_vector(to_unsigned(6295, LDPC_TABLE_DATA_WIDTH)),
    2312 => std_logic_vector(to_unsigned(11329, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2313 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    2314 => std_logic_vector(to_unsigned(1409, LDPC_TABLE_DATA_WIDTH)),
    2315 => std_logic_vector(to_unsigned(12061, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2316 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    2317 => std_logic_vector(to_unsigned(8065, LDPC_TABLE_DATA_WIDTH)),
    2318 => std_logic_vector(to_unsigned(9087, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2319 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    2320 => std_logic_vector(to_unsigned(2918, LDPC_TABLE_DATA_WIDTH)),
    2321 => std_logic_vector(to_unsigned(8438, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2322 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    2323 => std_logic_vector(to_unsigned(1293, LDPC_TABLE_DATA_WIDTH)),
    2324 => std_logic_vector(to_unsigned(14115, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2325 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    2326 => std_logic_vector(to_unsigned(3922, LDPC_TABLE_DATA_WIDTH)),
    2327 => std_logic_vector(to_unsigned(13851, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2328 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    2329 => std_logic_vector(to_unsigned(3851, LDPC_TABLE_DATA_WIDTH)),
    2330 => std_logic_vector(to_unsigned(4000, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2331 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    2332 => std_logic_vector(to_unsigned(5865, LDPC_TABLE_DATA_WIDTH)),
    2333 => std_logic_vector(to_unsigned(1768, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2334 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    2335 => std_logic_vector(to_unsigned(2655, LDPC_TABLE_DATA_WIDTH)),
    2336 => std_logic_vector(to_unsigned(14957, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2337 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    2338 => std_logic_vector(to_unsigned(5565, LDPC_TABLE_DATA_WIDTH)),
    2339 => std_logic_vector(to_unsigned(6332, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2340 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    2341 => std_logic_vector(to_unsigned(4303, LDPC_TABLE_DATA_WIDTH)),
    2342 => std_logic_vector(to_unsigned(12631, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2343 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    2344 => std_logic_vector(to_unsigned(11653, LDPC_TABLE_DATA_WIDTH)),
    2345 => std_logic_vector(to_unsigned(12236, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2346 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    2347 => std_logic_vector(to_unsigned(16025, LDPC_TABLE_DATA_WIDTH)),
    2348 => std_logic_vector(to_unsigned(7632, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2349 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    2350 => std_logic_vector(to_unsigned(4655, LDPC_TABLE_DATA_WIDTH)),
    2351 => std_logic_vector(to_unsigned(14128, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2352 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    2353 => std_logic_vector(to_unsigned(9584, LDPC_TABLE_DATA_WIDTH)),
    2354 => std_logic_vector(to_unsigned(13123, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2355 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    2356 => std_logic_vector(to_unsigned(13987, LDPC_TABLE_DATA_WIDTH)),
    2357 => std_logic_vector(to_unsigned(9597, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2358 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    2359 => std_logic_vector(to_unsigned(15409, LDPC_TABLE_DATA_WIDTH)),
    2360 => std_logic_vector(to_unsigned(12110, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2361 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    2362 => std_logic_vector(to_unsigned(8754, LDPC_TABLE_DATA_WIDTH)),
    2363 => std_logic_vector(to_unsigned(15490, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2364 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    2365 => std_logic_vector(to_unsigned(7416, LDPC_TABLE_DATA_WIDTH)),
    2366 => std_logic_vector(to_unsigned(15325, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2367 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    2368 => std_logic_vector(to_unsigned(2909, LDPC_TABLE_DATA_WIDTH)),
    2369 => std_logic_vector(to_unsigned(15549, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2370 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    2371 => std_logic_vector(to_unsigned(2995, LDPC_TABLE_DATA_WIDTH)),
    2372 => std_logic_vector(to_unsigned(8257, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2373 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    2374 => std_logic_vector(to_unsigned(9406, LDPC_TABLE_DATA_WIDTH)),
    2375 => std_logic_vector(to_unsigned(4791, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2376 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    2377 => std_logic_vector(to_unsigned(11111, LDPC_TABLE_DATA_WIDTH)),
    2378 => std_logic_vector(to_unsigned(4854, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2379 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    2380 => std_logic_vector(to_unsigned(2812, LDPC_TABLE_DATA_WIDTH)),
    2381 => std_logic_vector(to_unsigned(8521, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2382 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    2383 => std_logic_vector(to_unsigned(8476, LDPC_TABLE_DATA_WIDTH)),
    2384 => std_logic_vector(to_unsigned(14717, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2385 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    2386 => std_logic_vector(to_unsigned(7820, LDPC_TABLE_DATA_WIDTH)),
    2387 => std_logic_vector(to_unsigned(15360, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2388 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    2389 => std_logic_vector(to_unsigned(1179, LDPC_TABLE_DATA_WIDTH)),
    2390 => std_logic_vector(to_unsigned(7939, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2391 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    2392 => std_logic_vector(to_unsigned(2357, LDPC_TABLE_DATA_WIDTH)),
    2393 => std_logic_vector(to_unsigned(8678, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2394 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    2395 => std_logic_vector(to_unsigned(7703, LDPC_TABLE_DATA_WIDTH)),
    2396 => std_logic_vector(to_unsigned(6216, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2397 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    2398 => std_logic_vector(to_unsigned(3477, LDPC_TABLE_DATA_WIDTH)),
    2399 => std_logic_vector(to_unsigned(7067, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2400 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    2401 => std_logic_vector(to_unsigned(3931, LDPC_TABLE_DATA_WIDTH)),
    2402 => std_logic_vector(to_unsigned(13845, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2403 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    2404 => std_logic_vector(to_unsigned(7675, LDPC_TABLE_DATA_WIDTH)),
    2405 => std_logic_vector(to_unsigned(12899, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2406 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    2407 => std_logic_vector(to_unsigned(1754, LDPC_TABLE_DATA_WIDTH)),
    2408 => std_logic_vector(to_unsigned(8187, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2409 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    2410 => std_logic_vector(to_unsigned(7785, LDPC_TABLE_DATA_WIDTH)),
    2411 => std_logic_vector(to_unsigned(1400, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2412 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    2413 => std_logic_vector(to_unsigned(9213, LDPC_TABLE_DATA_WIDTH)),
    2414 => std_logic_vector(to_unsigned(5891, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2415 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    2416 => std_logic_vector(to_unsigned(2494, LDPC_TABLE_DATA_WIDTH)),
    2417 => std_logic_vector(to_unsigned(7703, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2418 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    2419 => std_logic_vector(to_unsigned(2576, LDPC_TABLE_DATA_WIDTH)),
    2420 => std_logic_vector(to_unsigned(7902, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2421 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    2422 => std_logic_vector(to_unsigned(4821, LDPC_TABLE_DATA_WIDTH)),
    2423 => std_logic_vector(to_unsigned(15682, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2424 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    2425 => std_logic_vector(to_unsigned(10426, LDPC_TABLE_DATA_WIDTH)),
    2426 => std_logic_vector(to_unsigned(11935, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2427 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    2428 => std_logic_vector(to_unsigned(1810, LDPC_TABLE_DATA_WIDTH)),
    2429 => std_logic_vector(to_unsigned(904, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2430 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    2431 => std_logic_vector(to_unsigned(11332, LDPC_TABLE_DATA_WIDTH)),
    2432 => std_logic_vector(to_unsigned(9264, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2433 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    2434 => std_logic_vector(to_unsigned(11312, LDPC_TABLE_DATA_WIDTH)),
    2435 => std_logic_vector(to_unsigned(3570, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2436 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    2437 => std_logic_vector(to_unsigned(14916, LDPC_TABLE_DATA_WIDTH)),
    2438 => std_logic_vector(to_unsigned(2650, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2439 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    2440 => std_logic_vector(to_unsigned(7679, LDPC_TABLE_DATA_WIDTH)),
    2441 => std_logic_vector(to_unsigned(7842, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2442 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    2443 => std_logic_vector(to_unsigned(6089, LDPC_TABLE_DATA_WIDTH)),
    2444 => std_logic_vector(to_unsigned(13084, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2445 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    2446 => std_logic_vector(to_unsigned(3938, LDPC_TABLE_DATA_WIDTH)),
    2447 => std_logic_vector(to_unsigned(2751, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2448 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    2449 => std_logic_vector(to_unsigned(8509, LDPC_TABLE_DATA_WIDTH)),
    2450 => std_logic_vector(to_unsigned(4648, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2451 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    2452 => std_logic_vector(to_unsigned(12204, LDPC_TABLE_DATA_WIDTH)),
    2453 => std_logic_vector(to_unsigned(8917, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2454 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    2455 => std_logic_vector(to_unsigned(5749, LDPC_TABLE_DATA_WIDTH)),
    2456 => std_logic_vector(to_unsigned(12443, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2457 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    2458 => std_logic_vector(to_unsigned(12613, LDPC_TABLE_DATA_WIDTH)),
    2459 => std_logic_vector(to_unsigned(4431, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2460 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    2461 => std_logic_vector(to_unsigned(1344, LDPC_TABLE_DATA_WIDTH)),
    2462 => std_logic_vector(to_unsigned(4014, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2463 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    2464 => std_logic_vector(to_unsigned(8488, LDPC_TABLE_DATA_WIDTH)),
    2465 => std_logic_vector(to_unsigned(13850, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2466 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    2467 => std_logic_vector(to_unsigned(1730, LDPC_TABLE_DATA_WIDTH)),
    2468 => std_logic_vector(to_unsigned(14896, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2469 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    2470 => std_logic_vector(to_unsigned(14942, LDPC_TABLE_DATA_WIDTH)),
    2471 => std_logic_vector(to_unsigned(7126, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2472 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    2473 => std_logic_vector(to_unsigned(14983, LDPC_TABLE_DATA_WIDTH)),
    2474 => std_logic_vector(to_unsigned(8863, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2475 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    2476 => std_logic_vector(to_unsigned(6578, LDPC_TABLE_DATA_WIDTH)),
    2477 => std_logic_vector(to_unsigned(8564, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2478 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    2479 => std_logic_vector(to_unsigned(4947, LDPC_TABLE_DATA_WIDTH)),
    2480 => std_logic_vector(to_unsigned(396, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2481 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    2482 => std_logic_vector(to_unsigned(297, LDPC_TABLE_DATA_WIDTH)),
    2483 => std_logic_vector(to_unsigned(12805, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2484 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    2485 => std_logic_vector(to_unsigned(13878, LDPC_TABLE_DATA_WIDTH)),
    2486 => std_logic_vector(to_unsigned(6692, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2487 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    2488 => std_logic_vector(to_unsigned(11857, LDPC_TABLE_DATA_WIDTH)),
    2489 => std_logic_vector(to_unsigned(11186, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2490 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    2491 => std_logic_vector(to_unsigned(14395, LDPC_TABLE_DATA_WIDTH)),
    2492 => std_logic_vector(to_unsigned(11493, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2493 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    2494 => std_logic_vector(to_unsigned(16145, LDPC_TABLE_DATA_WIDTH)),
    2495 => std_logic_vector(to_unsigned(12251, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2496 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    2497 => std_logic_vector(to_unsigned(13462, LDPC_TABLE_DATA_WIDTH)),
    2498 => std_logic_vector(to_unsigned(7428, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2499 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    2500 => std_logic_vector(to_unsigned(14526, LDPC_TABLE_DATA_WIDTH)),
    2501 => std_logic_vector(to_unsigned(13119, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2502 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    2503 => std_logic_vector(to_unsigned(2535, LDPC_TABLE_DATA_WIDTH)),
    2504 => std_logic_vector(to_unsigned(11243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2505 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    2506 => std_logic_vector(to_unsigned(6465, LDPC_TABLE_DATA_WIDTH)),
    2507 => std_logic_vector(to_unsigned(12690, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2508 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    2509 => std_logic_vector(to_unsigned(6872, LDPC_TABLE_DATA_WIDTH)),
    2510 => std_logic_vector(to_unsigned(9334, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2511 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    2512 => std_logic_vector(to_unsigned(15371, LDPC_TABLE_DATA_WIDTH)),
    2513 => std_logic_vector(to_unsigned(14023, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2514 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    2515 => std_logic_vector(to_unsigned(8101, LDPC_TABLE_DATA_WIDTH)),
    2516 => std_logic_vector(to_unsigned(10187, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2517 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    2518 => std_logic_vector(to_unsigned(11963, LDPC_TABLE_DATA_WIDTH)),
    2519 => std_logic_vector(to_unsigned(4848, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2520 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    2521 => std_logic_vector(to_unsigned(15125, LDPC_TABLE_DATA_WIDTH)),
    2522 => std_logic_vector(to_unsigned(6119, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2523 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    2524 => std_logic_vector(to_unsigned(8051, LDPC_TABLE_DATA_WIDTH)),
    2525 => std_logic_vector(to_unsigned(14465, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2526 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    2527 => std_logic_vector(to_unsigned(11139, LDPC_TABLE_DATA_WIDTH)),
    2528 => std_logic_vector(to_unsigned(5167, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2529 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    2530 => std_logic_vector(to_unsigned(2883, LDPC_TABLE_DATA_WIDTH)),
    2531 => std_logic_vector(to_unsigned(14521, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C3_5
    2532 => std_logic_vector(to_unsigned(22422, LDPC_TABLE_DATA_WIDTH)),
    2533 => std_logic_vector(to_unsigned(10282, LDPC_TABLE_DATA_WIDTH)),
    2534 => std_logic_vector(to_unsigned(11626, LDPC_TABLE_DATA_WIDTH)),
    2535 => std_logic_vector(to_unsigned(19997, LDPC_TABLE_DATA_WIDTH)),
    2536 => std_logic_vector(to_unsigned(11161, LDPC_TABLE_DATA_WIDTH)),
    2537 => std_logic_vector(to_unsigned(2922, LDPC_TABLE_DATA_WIDTH)),
    2538 => std_logic_vector(to_unsigned(3122, LDPC_TABLE_DATA_WIDTH)),
    2539 => std_logic_vector(to_unsigned(99, LDPC_TABLE_DATA_WIDTH)),
    2540 => std_logic_vector(to_unsigned(5625, LDPC_TABLE_DATA_WIDTH)),
    2541 => std_logic_vector(to_unsigned(17064, LDPC_TABLE_DATA_WIDTH)),
    2542 => std_logic_vector(to_unsigned(8270, LDPC_TABLE_DATA_WIDTH)),
    2543 => std_logic_vector(to_unsigned(179, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2544 => std_logic_vector(to_unsigned(25087, LDPC_TABLE_DATA_WIDTH)),
    2545 => std_logic_vector(to_unsigned(16218, LDPC_TABLE_DATA_WIDTH)),
    2546 => std_logic_vector(to_unsigned(17015, LDPC_TABLE_DATA_WIDTH)),
    2547 => std_logic_vector(to_unsigned(828, LDPC_TABLE_DATA_WIDTH)),
    2548 => std_logic_vector(to_unsigned(20041, LDPC_TABLE_DATA_WIDTH)),
    2549 => std_logic_vector(to_unsigned(25656, LDPC_TABLE_DATA_WIDTH)),
    2550 => std_logic_vector(to_unsigned(4186, LDPC_TABLE_DATA_WIDTH)),
    2551 => std_logic_vector(to_unsigned(11629, LDPC_TABLE_DATA_WIDTH)),
    2552 => std_logic_vector(to_unsigned(22599, LDPC_TABLE_DATA_WIDTH)),
    2553 => std_logic_vector(to_unsigned(17305, LDPC_TABLE_DATA_WIDTH)),
    2554 => std_logic_vector(to_unsigned(22515, LDPC_TABLE_DATA_WIDTH)),
    2555 => std_logic_vector(to_unsigned(6463, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2556 => std_logic_vector(to_unsigned(11049, LDPC_TABLE_DATA_WIDTH)),
    2557 => std_logic_vector(to_unsigned(22853, LDPC_TABLE_DATA_WIDTH)),
    2558 => std_logic_vector(to_unsigned(25706, LDPC_TABLE_DATA_WIDTH)),
    2559 => std_logic_vector(to_unsigned(14388, LDPC_TABLE_DATA_WIDTH)),
    2560 => std_logic_vector(to_unsigned(5500, LDPC_TABLE_DATA_WIDTH)),
    2561 => std_logic_vector(to_unsigned(19245, LDPC_TABLE_DATA_WIDTH)),
    2562 => std_logic_vector(to_unsigned(8732, LDPC_TABLE_DATA_WIDTH)),
    2563 => std_logic_vector(to_unsigned(2177, LDPC_TABLE_DATA_WIDTH)),
    2564 => std_logic_vector(to_unsigned(13555, LDPC_TABLE_DATA_WIDTH)),
    2565 => std_logic_vector(to_unsigned(11346, LDPC_TABLE_DATA_WIDTH)),
    2566 => std_logic_vector(to_unsigned(17265, LDPC_TABLE_DATA_WIDTH)),
    2567 => std_logic_vector(to_unsigned(3069, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2568 => std_logic_vector(to_unsigned(16581, LDPC_TABLE_DATA_WIDTH)),
    2569 => std_logic_vector(to_unsigned(22225, LDPC_TABLE_DATA_WIDTH)),
    2570 => std_logic_vector(to_unsigned(12563, LDPC_TABLE_DATA_WIDTH)),
    2571 => std_logic_vector(to_unsigned(19717, LDPC_TABLE_DATA_WIDTH)),
    2572 => std_logic_vector(to_unsigned(23577, LDPC_TABLE_DATA_WIDTH)),
    2573 => std_logic_vector(to_unsigned(11555, LDPC_TABLE_DATA_WIDTH)),
    2574 => std_logic_vector(to_unsigned(25496, LDPC_TABLE_DATA_WIDTH)),
    2575 => std_logic_vector(to_unsigned(6853, LDPC_TABLE_DATA_WIDTH)),
    2576 => std_logic_vector(to_unsigned(25403, LDPC_TABLE_DATA_WIDTH)),
    2577 => std_logic_vector(to_unsigned(5218, LDPC_TABLE_DATA_WIDTH)),
    2578 => std_logic_vector(to_unsigned(15925, LDPC_TABLE_DATA_WIDTH)),
    2579 => std_logic_vector(to_unsigned(21766, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2580 => std_logic_vector(to_unsigned(16529, LDPC_TABLE_DATA_WIDTH)),
    2581 => std_logic_vector(to_unsigned(14487, LDPC_TABLE_DATA_WIDTH)),
    2582 => std_logic_vector(to_unsigned(7643, LDPC_TABLE_DATA_WIDTH)),
    2583 => std_logic_vector(to_unsigned(10715, LDPC_TABLE_DATA_WIDTH)),
    2584 => std_logic_vector(to_unsigned(17442, LDPC_TABLE_DATA_WIDTH)),
    2585 => std_logic_vector(to_unsigned(11119, LDPC_TABLE_DATA_WIDTH)),
    2586 => std_logic_vector(to_unsigned(5679, LDPC_TABLE_DATA_WIDTH)),
    2587 => std_logic_vector(to_unsigned(14155, LDPC_TABLE_DATA_WIDTH)),
    2588 => std_logic_vector(to_unsigned(24213, LDPC_TABLE_DATA_WIDTH)),
    2589 => std_logic_vector(to_unsigned(21000, LDPC_TABLE_DATA_WIDTH)),
    2590 => std_logic_vector(to_unsigned(1116, LDPC_TABLE_DATA_WIDTH)),
    2591 => std_logic_vector(to_unsigned(15620, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2592 => std_logic_vector(to_unsigned(5340, LDPC_TABLE_DATA_WIDTH)),
    2593 => std_logic_vector(to_unsigned(8636, LDPC_TABLE_DATA_WIDTH)),
    2594 => std_logic_vector(to_unsigned(16693, LDPC_TABLE_DATA_WIDTH)),
    2595 => std_logic_vector(to_unsigned(1434, LDPC_TABLE_DATA_WIDTH)),
    2596 => std_logic_vector(to_unsigned(5635, LDPC_TABLE_DATA_WIDTH)),
    2597 => std_logic_vector(to_unsigned(6516, LDPC_TABLE_DATA_WIDTH)),
    2598 => std_logic_vector(to_unsigned(9482, LDPC_TABLE_DATA_WIDTH)),
    2599 => std_logic_vector(to_unsigned(20189, LDPC_TABLE_DATA_WIDTH)),
    2600 => std_logic_vector(to_unsigned(1066, LDPC_TABLE_DATA_WIDTH)),
    2601 => std_logic_vector(to_unsigned(15013, LDPC_TABLE_DATA_WIDTH)),
    2602 => std_logic_vector(to_unsigned(25361, LDPC_TABLE_DATA_WIDTH)),
    2603 => std_logic_vector(to_unsigned(14243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2604 => std_logic_vector(to_unsigned(18506, LDPC_TABLE_DATA_WIDTH)),
    2605 => std_logic_vector(to_unsigned(22236, LDPC_TABLE_DATA_WIDTH)),
    2606 => std_logic_vector(to_unsigned(20912, LDPC_TABLE_DATA_WIDTH)),
    2607 => std_logic_vector(to_unsigned(8952, LDPC_TABLE_DATA_WIDTH)),
    2608 => std_logic_vector(to_unsigned(5421, LDPC_TABLE_DATA_WIDTH)),
    2609 => std_logic_vector(to_unsigned(15691, LDPC_TABLE_DATA_WIDTH)),
    2610 => std_logic_vector(to_unsigned(6126, LDPC_TABLE_DATA_WIDTH)),
    2611 => std_logic_vector(to_unsigned(21595, LDPC_TABLE_DATA_WIDTH)),
    2612 => std_logic_vector(to_unsigned(500, LDPC_TABLE_DATA_WIDTH)),
    2613 => std_logic_vector(to_unsigned(6904, LDPC_TABLE_DATA_WIDTH)),
    2614 => std_logic_vector(to_unsigned(13059, LDPC_TABLE_DATA_WIDTH)),
    2615 => std_logic_vector(to_unsigned(6802, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2616 => std_logic_vector(to_unsigned(8433, LDPC_TABLE_DATA_WIDTH)),
    2617 => std_logic_vector(to_unsigned(4694, LDPC_TABLE_DATA_WIDTH)),
    2618 => std_logic_vector(to_unsigned(5524, LDPC_TABLE_DATA_WIDTH)),
    2619 => std_logic_vector(to_unsigned(14216, LDPC_TABLE_DATA_WIDTH)),
    2620 => std_logic_vector(to_unsigned(3685, LDPC_TABLE_DATA_WIDTH)),
    2621 => std_logic_vector(to_unsigned(19721, LDPC_TABLE_DATA_WIDTH)),
    2622 => std_logic_vector(to_unsigned(25420, LDPC_TABLE_DATA_WIDTH)),
    2623 => std_logic_vector(to_unsigned(9937, LDPC_TABLE_DATA_WIDTH)),
    2624 => std_logic_vector(to_unsigned(23813, LDPC_TABLE_DATA_WIDTH)),
    2625 => std_logic_vector(to_unsigned(9047, LDPC_TABLE_DATA_WIDTH)),
    2626 => std_logic_vector(to_unsigned(25651, LDPC_TABLE_DATA_WIDTH)),
    2627 => std_logic_vector(to_unsigned(16826, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2628 => std_logic_vector(to_unsigned(21500, LDPC_TABLE_DATA_WIDTH)),
    2629 => std_logic_vector(to_unsigned(24814, LDPC_TABLE_DATA_WIDTH)),
    2630 => std_logic_vector(to_unsigned(6344, LDPC_TABLE_DATA_WIDTH)),
    2631 => std_logic_vector(to_unsigned(17382, LDPC_TABLE_DATA_WIDTH)),
    2632 => std_logic_vector(to_unsigned(7064, LDPC_TABLE_DATA_WIDTH)),
    2633 => std_logic_vector(to_unsigned(13929, LDPC_TABLE_DATA_WIDTH)),
    2634 => std_logic_vector(to_unsigned(4004, LDPC_TABLE_DATA_WIDTH)),
    2635 => std_logic_vector(to_unsigned(16552, LDPC_TABLE_DATA_WIDTH)),
    2636 => std_logic_vector(to_unsigned(12818, LDPC_TABLE_DATA_WIDTH)),
    2637 => std_logic_vector(to_unsigned(8720, LDPC_TABLE_DATA_WIDTH)),
    2638 => std_logic_vector(to_unsigned(5286, LDPC_TABLE_DATA_WIDTH)),
    2639 => std_logic_vector(to_unsigned(2206, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2640 => std_logic_vector(to_unsigned(22517, LDPC_TABLE_DATA_WIDTH)),
    2641 => std_logic_vector(to_unsigned(2429, LDPC_TABLE_DATA_WIDTH)),
    2642 => std_logic_vector(to_unsigned(19065, LDPC_TABLE_DATA_WIDTH)),
    2643 => std_logic_vector(to_unsigned(2921, LDPC_TABLE_DATA_WIDTH)),
    2644 => std_logic_vector(to_unsigned(21611, LDPC_TABLE_DATA_WIDTH)),
    2645 => std_logic_vector(to_unsigned(1873, LDPC_TABLE_DATA_WIDTH)),
    2646 => std_logic_vector(to_unsigned(7507, LDPC_TABLE_DATA_WIDTH)),
    2647 => std_logic_vector(to_unsigned(5661, LDPC_TABLE_DATA_WIDTH)),
    2648 => std_logic_vector(to_unsigned(23006, LDPC_TABLE_DATA_WIDTH)),
    2649 => std_logic_vector(to_unsigned(23128, LDPC_TABLE_DATA_WIDTH)),
    2650 => std_logic_vector(to_unsigned(20543, LDPC_TABLE_DATA_WIDTH)),
    2651 => std_logic_vector(to_unsigned(19777, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2652 => std_logic_vector(to_unsigned(1770, LDPC_TABLE_DATA_WIDTH)),
    2653 => std_logic_vector(to_unsigned(4636, LDPC_TABLE_DATA_WIDTH)),
    2654 => std_logic_vector(to_unsigned(20900, LDPC_TABLE_DATA_WIDTH)),
    2655 => std_logic_vector(to_unsigned(14931, LDPC_TABLE_DATA_WIDTH)),
    2656 => std_logic_vector(to_unsigned(9247, LDPC_TABLE_DATA_WIDTH)),
    2657 => std_logic_vector(to_unsigned(12340, LDPC_TABLE_DATA_WIDTH)),
    2658 => std_logic_vector(to_unsigned(11008, LDPC_TABLE_DATA_WIDTH)),
    2659 => std_logic_vector(to_unsigned(12966, LDPC_TABLE_DATA_WIDTH)),
    2660 => std_logic_vector(to_unsigned(4471, LDPC_TABLE_DATA_WIDTH)),
    2661 => std_logic_vector(to_unsigned(2731, LDPC_TABLE_DATA_WIDTH)),
    2662 => std_logic_vector(to_unsigned(16445, LDPC_TABLE_DATA_WIDTH)),
    2663 => std_logic_vector(to_unsigned(791, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2664 => std_logic_vector(to_unsigned(6635, LDPC_TABLE_DATA_WIDTH)),
    2665 => std_logic_vector(to_unsigned(14556, LDPC_TABLE_DATA_WIDTH)),
    2666 => std_logic_vector(to_unsigned(18865, LDPC_TABLE_DATA_WIDTH)),
    2667 => std_logic_vector(to_unsigned(22421, LDPC_TABLE_DATA_WIDTH)),
    2668 => std_logic_vector(to_unsigned(22124, LDPC_TABLE_DATA_WIDTH)),
    2669 => std_logic_vector(to_unsigned(12697, LDPC_TABLE_DATA_WIDTH)),
    2670 => std_logic_vector(to_unsigned(9803, LDPC_TABLE_DATA_WIDTH)),
    2671 => std_logic_vector(to_unsigned(25485, LDPC_TABLE_DATA_WIDTH)),
    2672 => std_logic_vector(to_unsigned(7744, LDPC_TABLE_DATA_WIDTH)),
    2673 => std_logic_vector(to_unsigned(18254, LDPC_TABLE_DATA_WIDTH)),
    2674 => std_logic_vector(to_unsigned(11313, LDPC_TABLE_DATA_WIDTH)),
    2675 => std_logic_vector(to_unsigned(9004, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2676 => std_logic_vector(to_unsigned(19982, LDPC_TABLE_DATA_WIDTH)),
    2677 => std_logic_vector(to_unsigned(23963, LDPC_TABLE_DATA_WIDTH)),
    2678 => std_logic_vector(to_unsigned(18912, LDPC_TABLE_DATA_WIDTH)),
    2679 => std_logic_vector(to_unsigned(7206, LDPC_TABLE_DATA_WIDTH)),
    2680 => std_logic_vector(to_unsigned(12500, LDPC_TABLE_DATA_WIDTH)),
    2681 => std_logic_vector(to_unsigned(4382, LDPC_TABLE_DATA_WIDTH)),
    2682 => std_logic_vector(to_unsigned(20067, LDPC_TABLE_DATA_WIDTH)),
    2683 => std_logic_vector(to_unsigned(6177, LDPC_TABLE_DATA_WIDTH)),
    2684 => std_logic_vector(to_unsigned(21007, LDPC_TABLE_DATA_WIDTH)),
    2685 => std_logic_vector(to_unsigned(1195, LDPC_TABLE_DATA_WIDTH)),
    2686 => std_logic_vector(to_unsigned(23547, LDPC_TABLE_DATA_WIDTH)),
    2687 => std_logic_vector(to_unsigned(24837, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2688 => std_logic_vector(to_unsigned(756, LDPC_TABLE_DATA_WIDTH)),
    2689 => std_logic_vector(to_unsigned(11158, LDPC_TABLE_DATA_WIDTH)),
    2690 => std_logic_vector(to_unsigned(14646, LDPC_TABLE_DATA_WIDTH)),
    2691 => std_logic_vector(to_unsigned(20534, LDPC_TABLE_DATA_WIDTH)),
    2692 => std_logic_vector(to_unsigned(3647, LDPC_TABLE_DATA_WIDTH)),
    2693 => std_logic_vector(to_unsigned(17728, LDPC_TABLE_DATA_WIDTH)),
    2694 => std_logic_vector(to_unsigned(11676, LDPC_TABLE_DATA_WIDTH)),
    2695 => std_logic_vector(to_unsigned(11843, LDPC_TABLE_DATA_WIDTH)),
    2696 => std_logic_vector(to_unsigned(12937, LDPC_TABLE_DATA_WIDTH)),
    2697 => std_logic_vector(to_unsigned(4402, LDPC_TABLE_DATA_WIDTH)),
    2698 => std_logic_vector(to_unsigned(8261, LDPC_TABLE_DATA_WIDTH)),
    2699 => std_logic_vector(to_unsigned(22944, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2700 => std_logic_vector(to_unsigned(9306, LDPC_TABLE_DATA_WIDTH)),
    2701 => std_logic_vector(to_unsigned(24009, LDPC_TABLE_DATA_WIDTH)),
    2702 => std_logic_vector(to_unsigned(10012, LDPC_TABLE_DATA_WIDTH)),
    2703 => std_logic_vector(to_unsigned(11081, LDPC_TABLE_DATA_WIDTH)),
    2704 => std_logic_vector(to_unsigned(3746, LDPC_TABLE_DATA_WIDTH)),
    2705 => std_logic_vector(to_unsigned(24325, LDPC_TABLE_DATA_WIDTH)),
    2706 => std_logic_vector(to_unsigned(8060, LDPC_TABLE_DATA_WIDTH)),
    2707 => std_logic_vector(to_unsigned(19826, LDPC_TABLE_DATA_WIDTH)),
    2708 => std_logic_vector(to_unsigned(842, LDPC_TABLE_DATA_WIDTH)),
    2709 => std_logic_vector(to_unsigned(8836, LDPC_TABLE_DATA_WIDTH)),
    2710 => std_logic_vector(to_unsigned(2898, LDPC_TABLE_DATA_WIDTH)),
    2711 => std_logic_vector(to_unsigned(5019, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2712 => std_logic_vector(to_unsigned(7575, LDPC_TABLE_DATA_WIDTH)),
    2713 => std_logic_vector(to_unsigned(7455, LDPC_TABLE_DATA_WIDTH)),
    2714 => std_logic_vector(to_unsigned(25244, LDPC_TABLE_DATA_WIDTH)),
    2715 => std_logic_vector(to_unsigned(4736, LDPC_TABLE_DATA_WIDTH)),
    2716 => std_logic_vector(to_unsigned(14400, LDPC_TABLE_DATA_WIDTH)),
    2717 => std_logic_vector(to_unsigned(22981, LDPC_TABLE_DATA_WIDTH)),
    2718 => std_logic_vector(to_unsigned(5543, LDPC_TABLE_DATA_WIDTH)),
    2719 => std_logic_vector(to_unsigned(8006, LDPC_TABLE_DATA_WIDTH)),
    2720 => std_logic_vector(to_unsigned(24203, LDPC_TABLE_DATA_WIDTH)),
    2721 => std_logic_vector(to_unsigned(13053, LDPC_TABLE_DATA_WIDTH)),
    2722 => std_logic_vector(to_unsigned(1120, LDPC_TABLE_DATA_WIDTH)),
    2723 => std_logic_vector(to_unsigned(5128, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2724 => std_logic_vector(to_unsigned(3482, LDPC_TABLE_DATA_WIDTH)),
    2725 => std_logic_vector(to_unsigned(9270, LDPC_TABLE_DATA_WIDTH)),
    2726 => std_logic_vector(to_unsigned(13059, LDPC_TABLE_DATA_WIDTH)),
    2727 => std_logic_vector(to_unsigned(15825, LDPC_TABLE_DATA_WIDTH)),
    2728 => std_logic_vector(to_unsigned(7453, LDPC_TABLE_DATA_WIDTH)),
    2729 => std_logic_vector(to_unsigned(23747, LDPC_TABLE_DATA_WIDTH)),
    2730 => std_logic_vector(to_unsigned(3656, LDPC_TABLE_DATA_WIDTH)),
    2731 => std_logic_vector(to_unsigned(24585, LDPC_TABLE_DATA_WIDTH)),
    2732 => std_logic_vector(to_unsigned(16542, LDPC_TABLE_DATA_WIDTH)),
    2733 => std_logic_vector(to_unsigned(17507, LDPC_TABLE_DATA_WIDTH)),
    2734 => std_logic_vector(to_unsigned(22462, LDPC_TABLE_DATA_WIDTH)),
    2735 => std_logic_vector(to_unsigned(14670, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2736 => std_logic_vector(to_unsigned(15627, LDPC_TABLE_DATA_WIDTH)),
    2737 => std_logic_vector(to_unsigned(15290, LDPC_TABLE_DATA_WIDTH)),
    2738 => std_logic_vector(to_unsigned(4198, LDPC_TABLE_DATA_WIDTH)),
    2739 => std_logic_vector(to_unsigned(22748, LDPC_TABLE_DATA_WIDTH)),
    2740 => std_logic_vector(to_unsigned(5842, LDPC_TABLE_DATA_WIDTH)),
    2741 => std_logic_vector(to_unsigned(13395, LDPC_TABLE_DATA_WIDTH)),
    2742 => std_logic_vector(to_unsigned(23918, LDPC_TABLE_DATA_WIDTH)),
    2743 => std_logic_vector(to_unsigned(16985, LDPC_TABLE_DATA_WIDTH)),
    2744 => std_logic_vector(to_unsigned(14929, LDPC_TABLE_DATA_WIDTH)),
    2745 => std_logic_vector(to_unsigned(3726, LDPC_TABLE_DATA_WIDTH)),
    2746 => std_logic_vector(to_unsigned(25350, LDPC_TABLE_DATA_WIDTH)),
    2747 => std_logic_vector(to_unsigned(24157, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2748 => std_logic_vector(to_unsigned(24896, LDPC_TABLE_DATA_WIDTH)),
    2749 => std_logic_vector(to_unsigned(16365, LDPC_TABLE_DATA_WIDTH)),
    2750 => std_logic_vector(to_unsigned(16423, LDPC_TABLE_DATA_WIDTH)),
    2751 => std_logic_vector(to_unsigned(13461, LDPC_TABLE_DATA_WIDTH)),
    2752 => std_logic_vector(to_unsigned(16615, LDPC_TABLE_DATA_WIDTH)),
    2753 => std_logic_vector(to_unsigned(8107, LDPC_TABLE_DATA_WIDTH)),
    2754 => std_logic_vector(to_unsigned(24741, LDPC_TABLE_DATA_WIDTH)),
    2755 => std_logic_vector(to_unsigned(3604, LDPC_TABLE_DATA_WIDTH)),
    2756 => std_logic_vector(to_unsigned(25904, LDPC_TABLE_DATA_WIDTH)),
    2757 => std_logic_vector(to_unsigned(8716, LDPC_TABLE_DATA_WIDTH)),
    2758 => std_logic_vector(to_unsigned(9604, LDPC_TABLE_DATA_WIDTH)),
    2759 => std_logic_vector(to_unsigned(20365, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2760 => std_logic_vector(to_unsigned(3729, LDPC_TABLE_DATA_WIDTH)),
    2761 => std_logic_vector(to_unsigned(17245, LDPC_TABLE_DATA_WIDTH)),
    2762 => std_logic_vector(to_unsigned(18448, LDPC_TABLE_DATA_WIDTH)),
    2763 => std_logic_vector(to_unsigned(9862, LDPC_TABLE_DATA_WIDTH)),
    2764 => std_logic_vector(to_unsigned(20831, LDPC_TABLE_DATA_WIDTH)),
    2765 => std_logic_vector(to_unsigned(25326, LDPC_TABLE_DATA_WIDTH)),
    2766 => std_logic_vector(to_unsigned(20517, LDPC_TABLE_DATA_WIDTH)),
    2767 => std_logic_vector(to_unsigned(24618, LDPC_TABLE_DATA_WIDTH)),
    2768 => std_logic_vector(to_unsigned(13282, LDPC_TABLE_DATA_WIDTH)),
    2769 => std_logic_vector(to_unsigned(5099, LDPC_TABLE_DATA_WIDTH)),
    2770 => std_logic_vector(to_unsigned(14183, LDPC_TABLE_DATA_WIDTH)),
    2771 => std_logic_vector(to_unsigned(8804, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2772 => std_logic_vector(to_unsigned(16455, LDPC_TABLE_DATA_WIDTH)),
    2773 => std_logic_vector(to_unsigned(17646, LDPC_TABLE_DATA_WIDTH)),
    2774 => std_logic_vector(to_unsigned(15376, LDPC_TABLE_DATA_WIDTH)),
    2775 => std_logic_vector(to_unsigned(18194, LDPC_TABLE_DATA_WIDTH)),
    2776 => std_logic_vector(to_unsigned(25528, LDPC_TABLE_DATA_WIDTH)),
    2777 => std_logic_vector(to_unsigned(1777, LDPC_TABLE_DATA_WIDTH)),
    2778 => std_logic_vector(to_unsigned(6066, LDPC_TABLE_DATA_WIDTH)),
    2779 => std_logic_vector(to_unsigned(21855, LDPC_TABLE_DATA_WIDTH)),
    2780 => std_logic_vector(to_unsigned(14372, LDPC_TABLE_DATA_WIDTH)),
    2781 => std_logic_vector(to_unsigned(12517, LDPC_TABLE_DATA_WIDTH)),
    2782 => std_logic_vector(to_unsigned(4488, LDPC_TABLE_DATA_WIDTH)),
    2783 => std_logic_vector(to_unsigned(17490, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2784 => std_logic_vector(to_unsigned(1400, LDPC_TABLE_DATA_WIDTH)),
    2785 => std_logic_vector(to_unsigned(8135, LDPC_TABLE_DATA_WIDTH)),
    2786 => std_logic_vector(to_unsigned(23375, LDPC_TABLE_DATA_WIDTH)),
    2787 => std_logic_vector(to_unsigned(20879, LDPC_TABLE_DATA_WIDTH)),
    2788 => std_logic_vector(to_unsigned(8476, LDPC_TABLE_DATA_WIDTH)),
    2789 => std_logic_vector(to_unsigned(4084, LDPC_TABLE_DATA_WIDTH)),
    2790 => std_logic_vector(to_unsigned(12936, LDPC_TABLE_DATA_WIDTH)),
    2791 => std_logic_vector(to_unsigned(25536, LDPC_TABLE_DATA_WIDTH)),
    2792 => std_logic_vector(to_unsigned(22309, LDPC_TABLE_DATA_WIDTH)),
    2793 => std_logic_vector(to_unsigned(16582, LDPC_TABLE_DATA_WIDTH)),
    2794 => std_logic_vector(to_unsigned(6402, LDPC_TABLE_DATA_WIDTH)),
    2795 => std_logic_vector(to_unsigned(24360, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2796 => std_logic_vector(to_unsigned(25119, LDPC_TABLE_DATA_WIDTH)),
    2797 => std_logic_vector(to_unsigned(23586, LDPC_TABLE_DATA_WIDTH)),
    2798 => std_logic_vector(to_unsigned(128, LDPC_TABLE_DATA_WIDTH)),
    2799 => std_logic_vector(to_unsigned(4761, LDPC_TABLE_DATA_WIDTH)),
    2800 => std_logic_vector(to_unsigned(10443, LDPC_TABLE_DATA_WIDTH)),
    2801 => std_logic_vector(to_unsigned(22536, LDPC_TABLE_DATA_WIDTH)),
    2802 => std_logic_vector(to_unsigned(8607, LDPC_TABLE_DATA_WIDTH)),
    2803 => std_logic_vector(to_unsigned(9752, LDPC_TABLE_DATA_WIDTH)),
    2804 => std_logic_vector(to_unsigned(25446, LDPC_TABLE_DATA_WIDTH)),
    2805 => std_logic_vector(to_unsigned(15053, LDPC_TABLE_DATA_WIDTH)),
    2806 => std_logic_vector(to_unsigned(1856, LDPC_TABLE_DATA_WIDTH)),
    2807 => std_logic_vector(to_unsigned(4040, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2808 => std_logic_vector(to_unsigned(377, LDPC_TABLE_DATA_WIDTH)),
    2809 => std_logic_vector(to_unsigned(21160, LDPC_TABLE_DATA_WIDTH)),
    2810 => std_logic_vector(to_unsigned(13474, LDPC_TABLE_DATA_WIDTH)),
    2811 => std_logic_vector(to_unsigned(5451, LDPC_TABLE_DATA_WIDTH)),
    2812 => std_logic_vector(to_unsigned(17170, LDPC_TABLE_DATA_WIDTH)),
    2813 => std_logic_vector(to_unsigned(5938, LDPC_TABLE_DATA_WIDTH)),
    2814 => std_logic_vector(to_unsigned(10256, LDPC_TABLE_DATA_WIDTH)),
    2815 => std_logic_vector(to_unsigned(11972, LDPC_TABLE_DATA_WIDTH)),
    2816 => std_logic_vector(to_unsigned(24210, LDPC_TABLE_DATA_WIDTH)),
    2817 => std_logic_vector(to_unsigned(17833, LDPC_TABLE_DATA_WIDTH)),
    2818 => std_logic_vector(to_unsigned(22047, LDPC_TABLE_DATA_WIDTH)),
    2819 => std_logic_vector(to_unsigned(16108, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2820 => std_logic_vector(to_unsigned(13075, LDPC_TABLE_DATA_WIDTH)),
    2821 => std_logic_vector(to_unsigned(9648, LDPC_TABLE_DATA_WIDTH)),
    2822 => std_logic_vector(to_unsigned(24546, LDPC_TABLE_DATA_WIDTH)),
    2823 => std_logic_vector(to_unsigned(13150, LDPC_TABLE_DATA_WIDTH)),
    2824 => std_logic_vector(to_unsigned(23867, LDPC_TABLE_DATA_WIDTH)),
    2825 => std_logic_vector(to_unsigned(7309, LDPC_TABLE_DATA_WIDTH)),
    2826 => std_logic_vector(to_unsigned(19798, LDPC_TABLE_DATA_WIDTH)),
    2827 => std_logic_vector(to_unsigned(2988, LDPC_TABLE_DATA_WIDTH)),
    2828 => std_logic_vector(to_unsigned(16858, LDPC_TABLE_DATA_WIDTH)),
    2829 => std_logic_vector(to_unsigned(4825, LDPC_TABLE_DATA_WIDTH)),
    2830 => std_logic_vector(to_unsigned(23950, LDPC_TABLE_DATA_WIDTH)),
    2831 => std_logic_vector(to_unsigned(15125, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2832 => std_logic_vector(to_unsigned(20526, LDPC_TABLE_DATA_WIDTH)),
    2833 => std_logic_vector(to_unsigned(3553, LDPC_TABLE_DATA_WIDTH)),
    2834 => std_logic_vector(to_unsigned(11525, LDPC_TABLE_DATA_WIDTH)),
    2835 => std_logic_vector(to_unsigned(23366, LDPC_TABLE_DATA_WIDTH)),
    2836 => std_logic_vector(to_unsigned(2452, LDPC_TABLE_DATA_WIDTH)),
    2837 => std_logic_vector(to_unsigned(17626, LDPC_TABLE_DATA_WIDTH)),
    2838 => std_logic_vector(to_unsigned(19265, LDPC_TABLE_DATA_WIDTH)),
    2839 => std_logic_vector(to_unsigned(20172, LDPC_TABLE_DATA_WIDTH)),
    2840 => std_logic_vector(to_unsigned(18060, LDPC_TABLE_DATA_WIDTH)),
    2841 => std_logic_vector(to_unsigned(24593, LDPC_TABLE_DATA_WIDTH)),
    2842 => std_logic_vector(to_unsigned(13255, LDPC_TABLE_DATA_WIDTH)),
    2843 => std_logic_vector(to_unsigned(1552, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2844 => std_logic_vector(to_unsigned(18839, LDPC_TABLE_DATA_WIDTH)),
    2845 => std_logic_vector(to_unsigned(21132, LDPC_TABLE_DATA_WIDTH)),
    2846 => std_logic_vector(to_unsigned(20119, LDPC_TABLE_DATA_WIDTH)),
    2847 => std_logic_vector(to_unsigned(15214, LDPC_TABLE_DATA_WIDTH)),
    2848 => std_logic_vector(to_unsigned(14705, LDPC_TABLE_DATA_WIDTH)),
    2849 => std_logic_vector(to_unsigned(7096, LDPC_TABLE_DATA_WIDTH)),
    2850 => std_logic_vector(to_unsigned(10174, LDPC_TABLE_DATA_WIDTH)),
    2851 => std_logic_vector(to_unsigned(5663, LDPC_TABLE_DATA_WIDTH)),
    2852 => std_logic_vector(to_unsigned(18651, LDPC_TABLE_DATA_WIDTH)),
    2853 => std_logic_vector(to_unsigned(19700, LDPC_TABLE_DATA_WIDTH)),
    2854 => std_logic_vector(to_unsigned(12524, LDPC_TABLE_DATA_WIDTH)),
    2855 => std_logic_vector(to_unsigned(14033, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2856 => std_logic_vector(to_unsigned(4127, LDPC_TABLE_DATA_WIDTH)),
    2857 => std_logic_vector(to_unsigned(2971, LDPC_TABLE_DATA_WIDTH)),
    2858 => std_logic_vector(to_unsigned(17499, LDPC_TABLE_DATA_WIDTH)),
    2859 => std_logic_vector(to_unsigned(16287, LDPC_TABLE_DATA_WIDTH)),
    2860 => std_logic_vector(to_unsigned(22368, LDPC_TABLE_DATA_WIDTH)),
    2861 => std_logic_vector(to_unsigned(21463, LDPC_TABLE_DATA_WIDTH)),
    2862 => std_logic_vector(to_unsigned(7943, LDPC_TABLE_DATA_WIDTH)),
    2863 => std_logic_vector(to_unsigned(18880, LDPC_TABLE_DATA_WIDTH)),
    2864 => std_logic_vector(to_unsigned(5567, LDPC_TABLE_DATA_WIDTH)),
    2865 => std_logic_vector(to_unsigned(8047, LDPC_TABLE_DATA_WIDTH)),
    2866 => std_logic_vector(to_unsigned(23363, LDPC_TABLE_DATA_WIDTH)),
    2867 => std_logic_vector(to_unsigned(6797, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2868 => std_logic_vector(to_unsigned(10651, LDPC_TABLE_DATA_WIDTH)),
    2869 => std_logic_vector(to_unsigned(24471, LDPC_TABLE_DATA_WIDTH)),
    2870 => std_logic_vector(to_unsigned(14325, LDPC_TABLE_DATA_WIDTH)),
    2871 => std_logic_vector(to_unsigned(4081, LDPC_TABLE_DATA_WIDTH)),
    2872 => std_logic_vector(to_unsigned(7258, LDPC_TABLE_DATA_WIDTH)),
    2873 => std_logic_vector(to_unsigned(4949, LDPC_TABLE_DATA_WIDTH)),
    2874 => std_logic_vector(to_unsigned(7044, LDPC_TABLE_DATA_WIDTH)),
    2875 => std_logic_vector(to_unsigned(1078, LDPC_TABLE_DATA_WIDTH)),
    2876 => std_logic_vector(to_unsigned(797, LDPC_TABLE_DATA_WIDTH)),
    2877 => std_logic_vector(to_unsigned(22910, LDPC_TABLE_DATA_WIDTH)),
    2878 => std_logic_vector(to_unsigned(20474, LDPC_TABLE_DATA_WIDTH)),
    2879 => std_logic_vector(to_unsigned(4318, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2880 => std_logic_vector(to_unsigned(21374, LDPC_TABLE_DATA_WIDTH)),
    2881 => std_logic_vector(to_unsigned(13231, LDPC_TABLE_DATA_WIDTH)),
    2882 => std_logic_vector(to_unsigned(22985, LDPC_TABLE_DATA_WIDTH)),
    2883 => std_logic_vector(to_unsigned(5056, LDPC_TABLE_DATA_WIDTH)),
    2884 => std_logic_vector(to_unsigned(3821, LDPC_TABLE_DATA_WIDTH)),
    2885 => std_logic_vector(to_unsigned(23718, LDPC_TABLE_DATA_WIDTH)),
    2886 => std_logic_vector(to_unsigned(14178, LDPC_TABLE_DATA_WIDTH)),
    2887 => std_logic_vector(to_unsigned(9978, LDPC_TABLE_DATA_WIDTH)),
    2888 => std_logic_vector(to_unsigned(19030, LDPC_TABLE_DATA_WIDTH)),
    2889 => std_logic_vector(to_unsigned(23594, LDPC_TABLE_DATA_WIDTH)),
    2890 => std_logic_vector(to_unsigned(8895, LDPC_TABLE_DATA_WIDTH)),
    2891 => std_logic_vector(to_unsigned(25358, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2892 => std_logic_vector(to_unsigned(6199, LDPC_TABLE_DATA_WIDTH)),
    2893 => std_logic_vector(to_unsigned(22056, LDPC_TABLE_DATA_WIDTH)),
    2894 => std_logic_vector(to_unsigned(7749, LDPC_TABLE_DATA_WIDTH)),
    2895 => std_logic_vector(to_unsigned(13310, LDPC_TABLE_DATA_WIDTH)),
    2896 => std_logic_vector(to_unsigned(3999, LDPC_TABLE_DATA_WIDTH)),
    2897 => std_logic_vector(to_unsigned(23697, LDPC_TABLE_DATA_WIDTH)),
    2898 => std_logic_vector(to_unsigned(16445, LDPC_TABLE_DATA_WIDTH)),
    2899 => std_logic_vector(to_unsigned(22636, LDPC_TABLE_DATA_WIDTH)),
    2900 => std_logic_vector(to_unsigned(5225, LDPC_TABLE_DATA_WIDTH)),
    2901 => std_logic_vector(to_unsigned(22437, LDPC_TABLE_DATA_WIDTH)),
    2902 => std_logic_vector(to_unsigned(24153, LDPC_TABLE_DATA_WIDTH)),
    2903 => std_logic_vector(to_unsigned(9442, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2904 => std_logic_vector(to_unsigned(7978, LDPC_TABLE_DATA_WIDTH)),
    2905 => std_logic_vector(to_unsigned(12177, LDPC_TABLE_DATA_WIDTH)),
    2906 => std_logic_vector(to_unsigned(2893, LDPC_TABLE_DATA_WIDTH)),
    2907 => std_logic_vector(to_unsigned(20778, LDPC_TABLE_DATA_WIDTH)),
    2908 => std_logic_vector(to_unsigned(3175, LDPC_TABLE_DATA_WIDTH)),
    2909 => std_logic_vector(to_unsigned(8645, LDPC_TABLE_DATA_WIDTH)),
    2910 => std_logic_vector(to_unsigned(11863, LDPC_TABLE_DATA_WIDTH)),
    2911 => std_logic_vector(to_unsigned(24623, LDPC_TABLE_DATA_WIDTH)),
    2912 => std_logic_vector(to_unsigned(10311, LDPC_TABLE_DATA_WIDTH)),
    2913 => std_logic_vector(to_unsigned(25767, LDPC_TABLE_DATA_WIDTH)),
    2914 => std_logic_vector(to_unsigned(17057, LDPC_TABLE_DATA_WIDTH)),
    2915 => std_logic_vector(to_unsigned(3691, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2916 => std_logic_vector(to_unsigned(20473, LDPC_TABLE_DATA_WIDTH)),
    2917 => std_logic_vector(to_unsigned(11294, LDPC_TABLE_DATA_WIDTH)),
    2918 => std_logic_vector(to_unsigned(9914, LDPC_TABLE_DATA_WIDTH)),
    2919 => std_logic_vector(to_unsigned(22815, LDPC_TABLE_DATA_WIDTH)),
    2920 => std_logic_vector(to_unsigned(2574, LDPC_TABLE_DATA_WIDTH)),
    2921 => std_logic_vector(to_unsigned(8439, LDPC_TABLE_DATA_WIDTH)),
    2922 => std_logic_vector(to_unsigned(3699, LDPC_TABLE_DATA_WIDTH)),
    2923 => std_logic_vector(to_unsigned(5431, LDPC_TABLE_DATA_WIDTH)),
    2924 => std_logic_vector(to_unsigned(24840, LDPC_TABLE_DATA_WIDTH)),
    2925 => std_logic_vector(to_unsigned(21908, LDPC_TABLE_DATA_WIDTH)),
    2926 => std_logic_vector(to_unsigned(16088, LDPC_TABLE_DATA_WIDTH)),
    2927 => std_logic_vector(to_unsigned(18244, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2928 => std_logic_vector(to_unsigned(8208, LDPC_TABLE_DATA_WIDTH)),
    2929 => std_logic_vector(to_unsigned(5755, LDPC_TABLE_DATA_WIDTH)),
    2930 => std_logic_vector(to_unsigned(19059, LDPC_TABLE_DATA_WIDTH)),
    2931 => std_logic_vector(to_unsigned(8541, LDPC_TABLE_DATA_WIDTH)),
    2932 => std_logic_vector(to_unsigned(24924, LDPC_TABLE_DATA_WIDTH)),
    2933 => std_logic_vector(to_unsigned(6454, LDPC_TABLE_DATA_WIDTH)),
    2934 => std_logic_vector(to_unsigned(11234, LDPC_TABLE_DATA_WIDTH)),
    2935 => std_logic_vector(to_unsigned(10492, LDPC_TABLE_DATA_WIDTH)),
    2936 => std_logic_vector(to_unsigned(16406, LDPC_TABLE_DATA_WIDTH)),
    2937 => std_logic_vector(to_unsigned(10831, LDPC_TABLE_DATA_WIDTH)),
    2938 => std_logic_vector(to_unsigned(11436, LDPC_TABLE_DATA_WIDTH)),
    2939 => std_logic_vector(to_unsigned(9649, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2940 => std_logic_vector(to_unsigned(16264, LDPC_TABLE_DATA_WIDTH)),
    2941 => std_logic_vector(to_unsigned(11275, LDPC_TABLE_DATA_WIDTH)),
    2942 => std_logic_vector(to_unsigned(24953, LDPC_TABLE_DATA_WIDTH)),
    2943 => std_logic_vector(to_unsigned(2347, LDPC_TABLE_DATA_WIDTH)),
    2944 => std_logic_vector(to_unsigned(12667, LDPC_TABLE_DATA_WIDTH)),
    2945 => std_logic_vector(to_unsigned(19190, LDPC_TABLE_DATA_WIDTH)),
    2946 => std_logic_vector(to_unsigned(7257, LDPC_TABLE_DATA_WIDTH)),
    2947 => std_logic_vector(to_unsigned(7174, LDPC_TABLE_DATA_WIDTH)),
    2948 => std_logic_vector(to_unsigned(24819, LDPC_TABLE_DATA_WIDTH)),
    2949 => std_logic_vector(to_unsigned(2938, LDPC_TABLE_DATA_WIDTH)),
    2950 => std_logic_vector(to_unsigned(2522, LDPC_TABLE_DATA_WIDTH)),
    2951 => std_logic_vector(to_unsigned(11749, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2952 => std_logic_vector(to_unsigned(3627, LDPC_TABLE_DATA_WIDTH)),
    2953 => std_logic_vector(to_unsigned(5969, LDPC_TABLE_DATA_WIDTH)),
    2954 => std_logic_vector(to_unsigned(13862, LDPC_TABLE_DATA_WIDTH)),
    2955 => std_logic_vector(to_unsigned(1538, LDPC_TABLE_DATA_WIDTH)),
    2956 => std_logic_vector(to_unsigned(23176, LDPC_TABLE_DATA_WIDTH)),
    2957 => std_logic_vector(to_unsigned(6353, LDPC_TABLE_DATA_WIDTH)),
    2958 => std_logic_vector(to_unsigned(2855, LDPC_TABLE_DATA_WIDTH)),
    2959 => std_logic_vector(to_unsigned(17720, LDPC_TABLE_DATA_WIDTH)),
    2960 => std_logic_vector(to_unsigned(2472, LDPC_TABLE_DATA_WIDTH)),
    2961 => std_logic_vector(to_unsigned(7428, LDPC_TABLE_DATA_WIDTH)),
    2962 => std_logic_vector(to_unsigned(573, LDPC_TABLE_DATA_WIDTH)),
    2963 => std_logic_vector(to_unsigned(15036, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2964 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    2965 => std_logic_vector(to_unsigned(18539, LDPC_TABLE_DATA_WIDTH)),
    2966 => std_logic_vector(to_unsigned(18661, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2967 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    2968 => std_logic_vector(to_unsigned(10502, LDPC_TABLE_DATA_WIDTH)),
    2969 => std_logic_vector(to_unsigned(3002, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2970 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    2971 => std_logic_vector(to_unsigned(9368, LDPC_TABLE_DATA_WIDTH)),
    2972 => std_logic_vector(to_unsigned(10761, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2973 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    2974 => std_logic_vector(to_unsigned(12299, LDPC_TABLE_DATA_WIDTH)),
    2975 => std_logic_vector(to_unsigned(7828, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2976 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    2977 => std_logic_vector(to_unsigned(15048, LDPC_TABLE_DATA_WIDTH)),
    2978 => std_logic_vector(to_unsigned(13362, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2979 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    2980 => std_logic_vector(to_unsigned(18444, LDPC_TABLE_DATA_WIDTH)),
    2981 => std_logic_vector(to_unsigned(24640, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2982 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    2983 => std_logic_vector(to_unsigned(20775, LDPC_TABLE_DATA_WIDTH)),
    2984 => std_logic_vector(to_unsigned(19175, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2985 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    2986 => std_logic_vector(to_unsigned(18970, LDPC_TABLE_DATA_WIDTH)),
    2987 => std_logic_vector(to_unsigned(10971, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2988 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    2989 => std_logic_vector(to_unsigned(5329, LDPC_TABLE_DATA_WIDTH)),
    2990 => std_logic_vector(to_unsigned(19982, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2991 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    2992 => std_logic_vector(to_unsigned(11296, LDPC_TABLE_DATA_WIDTH)),
    2993 => std_logic_vector(to_unsigned(18655, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2994 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    2995 => std_logic_vector(to_unsigned(15046, LDPC_TABLE_DATA_WIDTH)),
    2996 => std_logic_vector(to_unsigned(20659, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    2997 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    2998 => std_logic_vector(to_unsigned(7300, LDPC_TABLE_DATA_WIDTH)),
    2999 => std_logic_vector(to_unsigned(22140, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3000 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3001 => std_logic_vector(to_unsigned(22029, LDPC_TABLE_DATA_WIDTH)),
    3002 => std_logic_vector(to_unsigned(14477, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3003 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3004 => std_logic_vector(to_unsigned(11129, LDPC_TABLE_DATA_WIDTH)),
    3005 => std_logic_vector(to_unsigned(742, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3006 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3007 => std_logic_vector(to_unsigned(13254, LDPC_TABLE_DATA_WIDTH)),
    3008 => std_logic_vector(to_unsigned(13813, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3009 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3010 => std_logic_vector(to_unsigned(19234, LDPC_TABLE_DATA_WIDTH)),
    3011 => std_logic_vector(to_unsigned(13273, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3012 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3013 => std_logic_vector(to_unsigned(6079, LDPC_TABLE_DATA_WIDTH)),
    3014 => std_logic_vector(to_unsigned(21122, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3015 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3016 => std_logic_vector(to_unsigned(22782, LDPC_TABLE_DATA_WIDTH)),
    3017 => std_logic_vector(to_unsigned(5828, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3018 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3019 => std_logic_vector(to_unsigned(19775, LDPC_TABLE_DATA_WIDTH)),
    3020 => std_logic_vector(to_unsigned(4247, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3021 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3022 => std_logic_vector(to_unsigned(1660, LDPC_TABLE_DATA_WIDTH)),
    3023 => std_logic_vector(to_unsigned(19413, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3024 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3025 => std_logic_vector(to_unsigned(4403, LDPC_TABLE_DATA_WIDTH)),
    3026 => std_logic_vector(to_unsigned(3649, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3027 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3028 => std_logic_vector(to_unsigned(13371, LDPC_TABLE_DATA_WIDTH)),
    3029 => std_logic_vector(to_unsigned(25851, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3030 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3031 => std_logic_vector(to_unsigned(22770, LDPC_TABLE_DATA_WIDTH)),
    3032 => std_logic_vector(to_unsigned(21784, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3033 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3034 => std_logic_vector(to_unsigned(10757, LDPC_TABLE_DATA_WIDTH)),
    3035 => std_logic_vector(to_unsigned(14131, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3036 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3037 => std_logic_vector(to_unsigned(16071, LDPC_TABLE_DATA_WIDTH)),
    3038 => std_logic_vector(to_unsigned(21617, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3039 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3040 => std_logic_vector(to_unsigned(6393, LDPC_TABLE_DATA_WIDTH)),
    3041 => std_logic_vector(to_unsigned(3725, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3042 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3043 => std_logic_vector(to_unsigned(597, LDPC_TABLE_DATA_WIDTH)),
    3044 => std_logic_vector(to_unsigned(19968, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3045 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3046 => std_logic_vector(to_unsigned(5743, LDPC_TABLE_DATA_WIDTH)),
    3047 => std_logic_vector(to_unsigned(8084, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3048 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3049 => std_logic_vector(to_unsigned(6770, LDPC_TABLE_DATA_WIDTH)),
    3050 => std_logic_vector(to_unsigned(9548, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3051 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3052 => std_logic_vector(to_unsigned(4285, LDPC_TABLE_DATA_WIDTH)),
    3053 => std_logic_vector(to_unsigned(17542, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3054 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    3055 => std_logic_vector(to_unsigned(13568, LDPC_TABLE_DATA_WIDTH)),
    3056 => std_logic_vector(to_unsigned(22599, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3057 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    3058 => std_logic_vector(to_unsigned(1786, LDPC_TABLE_DATA_WIDTH)),
    3059 => std_logic_vector(to_unsigned(4617, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3060 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    3061 => std_logic_vector(to_unsigned(23238, LDPC_TABLE_DATA_WIDTH)),
    3062 => std_logic_vector(to_unsigned(11648, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3063 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    3064 => std_logic_vector(to_unsigned(19627, LDPC_TABLE_DATA_WIDTH)),
    3065 => std_logic_vector(to_unsigned(2030, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3066 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    3067 => std_logic_vector(to_unsigned(13601, LDPC_TABLE_DATA_WIDTH)),
    3068 => std_logic_vector(to_unsigned(13458, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3069 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    3070 => std_logic_vector(to_unsigned(13740, LDPC_TABLE_DATA_WIDTH)),
    3071 => std_logic_vector(to_unsigned(17328, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3072 => std_logic_vector(to_unsigned(36, LDPC_TABLE_DATA_WIDTH)),
    3073 => std_logic_vector(to_unsigned(25012, LDPC_TABLE_DATA_WIDTH)),
    3074 => std_logic_vector(to_unsigned(13944, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3075 => std_logic_vector(to_unsigned(37, LDPC_TABLE_DATA_WIDTH)),
    3076 => std_logic_vector(to_unsigned(22513, LDPC_TABLE_DATA_WIDTH)),
    3077 => std_logic_vector(to_unsigned(6687, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3078 => std_logic_vector(to_unsigned(38, LDPC_TABLE_DATA_WIDTH)),
    3079 => std_logic_vector(to_unsigned(4934, LDPC_TABLE_DATA_WIDTH)),
    3080 => std_logic_vector(to_unsigned(12587, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3081 => std_logic_vector(to_unsigned(39, LDPC_TABLE_DATA_WIDTH)),
    3082 => std_logic_vector(to_unsigned(21197, LDPC_TABLE_DATA_WIDTH)),
    3083 => std_logic_vector(to_unsigned(5133, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3084 => std_logic_vector(to_unsigned(40, LDPC_TABLE_DATA_WIDTH)),
    3085 => std_logic_vector(to_unsigned(22705, LDPC_TABLE_DATA_WIDTH)),
    3086 => std_logic_vector(to_unsigned(6938, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3087 => std_logic_vector(to_unsigned(41, LDPC_TABLE_DATA_WIDTH)),
    3088 => std_logic_vector(to_unsigned(7534, LDPC_TABLE_DATA_WIDTH)),
    3089 => std_logic_vector(to_unsigned(24633, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3090 => std_logic_vector(to_unsigned(42, LDPC_TABLE_DATA_WIDTH)),
    3091 => std_logic_vector(to_unsigned(24400, LDPC_TABLE_DATA_WIDTH)),
    3092 => std_logic_vector(to_unsigned(12797, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3093 => std_logic_vector(to_unsigned(43, LDPC_TABLE_DATA_WIDTH)),
    3094 => std_logic_vector(to_unsigned(21911, LDPC_TABLE_DATA_WIDTH)),
    3095 => std_logic_vector(to_unsigned(25712, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3096 => std_logic_vector(to_unsigned(44, LDPC_TABLE_DATA_WIDTH)),
    3097 => std_logic_vector(to_unsigned(12039, LDPC_TABLE_DATA_WIDTH)),
    3098 => std_logic_vector(to_unsigned(1140, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3099 => std_logic_vector(to_unsigned(45, LDPC_TABLE_DATA_WIDTH)),
    3100 => std_logic_vector(to_unsigned(24306, LDPC_TABLE_DATA_WIDTH)),
    3101 => std_logic_vector(to_unsigned(1021, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3102 => std_logic_vector(to_unsigned(46, LDPC_TABLE_DATA_WIDTH)),
    3103 => std_logic_vector(to_unsigned(14012, LDPC_TABLE_DATA_WIDTH)),
    3104 => std_logic_vector(to_unsigned(20747, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3105 => std_logic_vector(to_unsigned(47, LDPC_TABLE_DATA_WIDTH)),
    3106 => std_logic_vector(to_unsigned(11265, LDPC_TABLE_DATA_WIDTH)),
    3107 => std_logic_vector(to_unsigned(15219, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3108 => std_logic_vector(to_unsigned(48, LDPC_TABLE_DATA_WIDTH)),
    3109 => std_logic_vector(to_unsigned(4670, LDPC_TABLE_DATA_WIDTH)),
    3110 => std_logic_vector(to_unsigned(15531, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3111 => std_logic_vector(to_unsigned(49, LDPC_TABLE_DATA_WIDTH)),
    3112 => std_logic_vector(to_unsigned(9417, LDPC_TABLE_DATA_WIDTH)),
    3113 => std_logic_vector(to_unsigned(14359, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3114 => std_logic_vector(to_unsigned(50, LDPC_TABLE_DATA_WIDTH)),
    3115 => std_logic_vector(to_unsigned(2415, LDPC_TABLE_DATA_WIDTH)),
    3116 => std_logic_vector(to_unsigned(6504, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3117 => std_logic_vector(to_unsigned(51, LDPC_TABLE_DATA_WIDTH)),
    3118 => std_logic_vector(to_unsigned(24964, LDPC_TABLE_DATA_WIDTH)),
    3119 => std_logic_vector(to_unsigned(24690, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3120 => std_logic_vector(to_unsigned(52, LDPC_TABLE_DATA_WIDTH)),
    3121 => std_logic_vector(to_unsigned(14443, LDPC_TABLE_DATA_WIDTH)),
    3122 => std_logic_vector(to_unsigned(8816, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3123 => std_logic_vector(to_unsigned(53, LDPC_TABLE_DATA_WIDTH)),
    3124 => std_logic_vector(to_unsigned(6926, LDPC_TABLE_DATA_WIDTH)),
    3125 => std_logic_vector(to_unsigned(1291, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3126 => std_logic_vector(to_unsigned(54, LDPC_TABLE_DATA_WIDTH)),
    3127 => std_logic_vector(to_unsigned(6209, LDPC_TABLE_DATA_WIDTH)),
    3128 => std_logic_vector(to_unsigned(20806, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3129 => std_logic_vector(to_unsigned(55, LDPC_TABLE_DATA_WIDTH)),
    3130 => std_logic_vector(to_unsigned(13915, LDPC_TABLE_DATA_WIDTH)),
    3131 => std_logic_vector(to_unsigned(4079, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3132 => std_logic_vector(to_unsigned(56, LDPC_TABLE_DATA_WIDTH)),
    3133 => std_logic_vector(to_unsigned(24410, LDPC_TABLE_DATA_WIDTH)),
    3134 => std_logic_vector(to_unsigned(13196, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3135 => std_logic_vector(to_unsigned(57, LDPC_TABLE_DATA_WIDTH)),
    3136 => std_logic_vector(to_unsigned(13505, LDPC_TABLE_DATA_WIDTH)),
    3137 => std_logic_vector(to_unsigned(6117, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3138 => std_logic_vector(to_unsigned(58, LDPC_TABLE_DATA_WIDTH)),
    3139 => std_logic_vector(to_unsigned(9869, LDPC_TABLE_DATA_WIDTH)),
    3140 => std_logic_vector(to_unsigned(8220, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3141 => std_logic_vector(to_unsigned(59, LDPC_TABLE_DATA_WIDTH)),
    3142 => std_logic_vector(to_unsigned(1570, LDPC_TABLE_DATA_WIDTH)),
    3143 => std_logic_vector(to_unsigned(6044, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3144 => std_logic_vector(to_unsigned(60, LDPC_TABLE_DATA_WIDTH)),
    3145 => std_logic_vector(to_unsigned(25780, LDPC_TABLE_DATA_WIDTH)),
    3146 => std_logic_vector(to_unsigned(17387, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3147 => std_logic_vector(to_unsigned(61, LDPC_TABLE_DATA_WIDTH)),
    3148 => std_logic_vector(to_unsigned(20671, LDPC_TABLE_DATA_WIDTH)),
    3149 => std_logic_vector(to_unsigned(24913, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3150 => std_logic_vector(to_unsigned(62, LDPC_TABLE_DATA_WIDTH)),
    3151 => std_logic_vector(to_unsigned(24558, LDPC_TABLE_DATA_WIDTH)),
    3152 => std_logic_vector(to_unsigned(20591, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3153 => std_logic_vector(to_unsigned(63, LDPC_TABLE_DATA_WIDTH)),
    3154 => std_logic_vector(to_unsigned(12402, LDPC_TABLE_DATA_WIDTH)),
    3155 => std_logic_vector(to_unsigned(3702, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3156 => std_logic_vector(to_unsigned(64, LDPC_TABLE_DATA_WIDTH)),
    3157 => std_logic_vector(to_unsigned(8314, LDPC_TABLE_DATA_WIDTH)),
    3158 => std_logic_vector(to_unsigned(1357, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3159 => std_logic_vector(to_unsigned(65, LDPC_TABLE_DATA_WIDTH)),
    3160 => std_logic_vector(to_unsigned(20071, LDPC_TABLE_DATA_WIDTH)),
    3161 => std_logic_vector(to_unsigned(14616, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3162 => std_logic_vector(to_unsigned(66, LDPC_TABLE_DATA_WIDTH)),
    3163 => std_logic_vector(to_unsigned(17014, LDPC_TABLE_DATA_WIDTH)),
    3164 => std_logic_vector(to_unsigned(3688, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3165 => std_logic_vector(to_unsigned(67, LDPC_TABLE_DATA_WIDTH)),
    3166 => std_logic_vector(to_unsigned(19837, LDPC_TABLE_DATA_WIDTH)),
    3167 => std_logic_vector(to_unsigned(946, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3168 => std_logic_vector(to_unsigned(68, LDPC_TABLE_DATA_WIDTH)),
    3169 => std_logic_vector(to_unsigned(15195, LDPC_TABLE_DATA_WIDTH)),
    3170 => std_logic_vector(to_unsigned(12136, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3171 => std_logic_vector(to_unsigned(69, LDPC_TABLE_DATA_WIDTH)),
    3172 => std_logic_vector(to_unsigned(7758, LDPC_TABLE_DATA_WIDTH)),
    3173 => std_logic_vector(to_unsigned(22808, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3174 => std_logic_vector(to_unsigned(70, LDPC_TABLE_DATA_WIDTH)),
    3175 => std_logic_vector(to_unsigned(3564, LDPC_TABLE_DATA_WIDTH)),
    3176 => std_logic_vector(to_unsigned(2925, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3177 => std_logic_vector(to_unsigned(71, LDPC_TABLE_DATA_WIDTH)),
    3178 => std_logic_vector(to_unsigned(3434, LDPC_TABLE_DATA_WIDTH)),
    3179 => std_logic_vector(to_unsigned(7769, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C4_5
    3180 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3181 => std_logic_vector(to_unsigned(149, LDPC_TABLE_DATA_WIDTH)),
    3182 => std_logic_vector(to_unsigned(11212, LDPC_TABLE_DATA_WIDTH)),
    3183 => std_logic_vector(to_unsigned(5575, LDPC_TABLE_DATA_WIDTH)),
    3184 => std_logic_vector(to_unsigned(6360, LDPC_TABLE_DATA_WIDTH)),
    3185 => std_logic_vector(to_unsigned(12559, LDPC_TABLE_DATA_WIDTH)),
    3186 => std_logic_vector(to_unsigned(8108, LDPC_TABLE_DATA_WIDTH)),
    3187 => std_logic_vector(to_unsigned(8505, LDPC_TABLE_DATA_WIDTH)),
    3188 => std_logic_vector(to_unsigned(408, LDPC_TABLE_DATA_WIDTH)),
    3189 => std_logic_vector(to_unsigned(10026, LDPC_TABLE_DATA_WIDTH)),
    3190 => std_logic_vector(to_unsigned(12828, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3191 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    3192 => std_logic_vector(to_unsigned(5237, LDPC_TABLE_DATA_WIDTH)),
    3193 => std_logic_vector(to_unsigned(490, LDPC_TABLE_DATA_WIDTH)),
    3194 => std_logic_vector(to_unsigned(10677, LDPC_TABLE_DATA_WIDTH)),
    3195 => std_logic_vector(to_unsigned(4998, LDPC_TABLE_DATA_WIDTH)),
    3196 => std_logic_vector(to_unsigned(3869, LDPC_TABLE_DATA_WIDTH)),
    3197 => std_logic_vector(to_unsigned(3734, LDPC_TABLE_DATA_WIDTH)),
    3198 => std_logic_vector(to_unsigned(3092, LDPC_TABLE_DATA_WIDTH)),
    3199 => std_logic_vector(to_unsigned(3509, LDPC_TABLE_DATA_WIDTH)),
    3200 => std_logic_vector(to_unsigned(7703, LDPC_TABLE_DATA_WIDTH)),
    3201 => std_logic_vector(to_unsigned(10305, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3202 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    3203 => std_logic_vector(to_unsigned(8742, LDPC_TABLE_DATA_WIDTH)),
    3204 => std_logic_vector(to_unsigned(5553, LDPC_TABLE_DATA_WIDTH)),
    3205 => std_logic_vector(to_unsigned(2820, LDPC_TABLE_DATA_WIDTH)),
    3206 => std_logic_vector(to_unsigned(7085, LDPC_TABLE_DATA_WIDTH)),
    3207 => std_logic_vector(to_unsigned(12116, LDPC_TABLE_DATA_WIDTH)),
    3208 => std_logic_vector(to_unsigned(10485, LDPC_TABLE_DATA_WIDTH)),
    3209 => std_logic_vector(to_unsigned(564, LDPC_TABLE_DATA_WIDTH)),
    3210 => std_logic_vector(to_unsigned(7795, LDPC_TABLE_DATA_WIDTH)),
    3211 => std_logic_vector(to_unsigned(2972, LDPC_TABLE_DATA_WIDTH)),
    3212 => std_logic_vector(to_unsigned(2157, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3213 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    3214 => std_logic_vector(to_unsigned(2699, LDPC_TABLE_DATA_WIDTH)),
    3215 => std_logic_vector(to_unsigned(4304, LDPC_TABLE_DATA_WIDTH)),
    3216 => std_logic_vector(to_unsigned(8350, LDPC_TABLE_DATA_WIDTH)),
    3217 => std_logic_vector(to_unsigned(712, LDPC_TABLE_DATA_WIDTH)),
    3218 => std_logic_vector(to_unsigned(2841, LDPC_TABLE_DATA_WIDTH)),
    3219 => std_logic_vector(to_unsigned(3250, LDPC_TABLE_DATA_WIDTH)),
    3220 => std_logic_vector(to_unsigned(4731, LDPC_TABLE_DATA_WIDTH)),
    3221 => std_logic_vector(to_unsigned(10105, LDPC_TABLE_DATA_WIDTH)),
    3222 => std_logic_vector(to_unsigned(517, LDPC_TABLE_DATA_WIDTH)),
    3223 => std_logic_vector(to_unsigned(7516, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3224 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    3225 => std_logic_vector(to_unsigned(12067, LDPC_TABLE_DATA_WIDTH)),
    3226 => std_logic_vector(to_unsigned(1351, LDPC_TABLE_DATA_WIDTH)),
    3227 => std_logic_vector(to_unsigned(11992, LDPC_TABLE_DATA_WIDTH)),
    3228 => std_logic_vector(to_unsigned(12191, LDPC_TABLE_DATA_WIDTH)),
    3229 => std_logic_vector(to_unsigned(11267, LDPC_TABLE_DATA_WIDTH)),
    3230 => std_logic_vector(to_unsigned(5161, LDPC_TABLE_DATA_WIDTH)),
    3231 => std_logic_vector(to_unsigned(537, LDPC_TABLE_DATA_WIDTH)),
    3232 => std_logic_vector(to_unsigned(6166, LDPC_TABLE_DATA_WIDTH)),
    3233 => std_logic_vector(to_unsigned(4246, LDPC_TABLE_DATA_WIDTH)),
    3234 => std_logic_vector(to_unsigned(2363, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3235 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    3236 => std_logic_vector(to_unsigned(6828, LDPC_TABLE_DATA_WIDTH)),
    3237 => std_logic_vector(to_unsigned(7107, LDPC_TABLE_DATA_WIDTH)),
    3238 => std_logic_vector(to_unsigned(2127, LDPC_TABLE_DATA_WIDTH)),
    3239 => std_logic_vector(to_unsigned(3724, LDPC_TABLE_DATA_WIDTH)),
    3240 => std_logic_vector(to_unsigned(5743, LDPC_TABLE_DATA_WIDTH)),
    3241 => std_logic_vector(to_unsigned(11040, LDPC_TABLE_DATA_WIDTH)),
    3242 => std_logic_vector(to_unsigned(10756, LDPC_TABLE_DATA_WIDTH)),
    3243 => std_logic_vector(to_unsigned(4073, LDPC_TABLE_DATA_WIDTH)),
    3244 => std_logic_vector(to_unsigned(1011, LDPC_TABLE_DATA_WIDTH)),
    3245 => std_logic_vector(to_unsigned(3422, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3246 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    3247 => std_logic_vector(to_unsigned(11259, LDPC_TABLE_DATA_WIDTH)),
    3248 => std_logic_vector(to_unsigned(1216, LDPC_TABLE_DATA_WIDTH)),
    3249 => std_logic_vector(to_unsigned(9526, LDPC_TABLE_DATA_WIDTH)),
    3250 => std_logic_vector(to_unsigned(1466, LDPC_TABLE_DATA_WIDTH)),
    3251 => std_logic_vector(to_unsigned(10816, LDPC_TABLE_DATA_WIDTH)),
    3252 => std_logic_vector(to_unsigned(940, LDPC_TABLE_DATA_WIDTH)),
    3253 => std_logic_vector(to_unsigned(3744, LDPC_TABLE_DATA_WIDTH)),
    3254 => std_logic_vector(to_unsigned(2815, LDPC_TABLE_DATA_WIDTH)),
    3255 => std_logic_vector(to_unsigned(11506, LDPC_TABLE_DATA_WIDTH)),
    3256 => std_logic_vector(to_unsigned(11573, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3257 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    3258 => std_logic_vector(to_unsigned(4549, LDPC_TABLE_DATA_WIDTH)),
    3259 => std_logic_vector(to_unsigned(11507, LDPC_TABLE_DATA_WIDTH)),
    3260 => std_logic_vector(to_unsigned(1118, LDPC_TABLE_DATA_WIDTH)),
    3261 => std_logic_vector(to_unsigned(1274, LDPC_TABLE_DATA_WIDTH)),
    3262 => std_logic_vector(to_unsigned(11751, LDPC_TABLE_DATA_WIDTH)),
    3263 => std_logic_vector(to_unsigned(5207, LDPC_TABLE_DATA_WIDTH)),
    3264 => std_logic_vector(to_unsigned(7854, LDPC_TABLE_DATA_WIDTH)),
    3265 => std_logic_vector(to_unsigned(12803, LDPC_TABLE_DATA_WIDTH)),
    3266 => std_logic_vector(to_unsigned(4047, LDPC_TABLE_DATA_WIDTH)),
    3267 => std_logic_vector(to_unsigned(6484, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3268 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    3269 => std_logic_vector(to_unsigned(8430, LDPC_TABLE_DATA_WIDTH)),
    3270 => std_logic_vector(to_unsigned(4115, LDPC_TABLE_DATA_WIDTH)),
    3271 => std_logic_vector(to_unsigned(9440, LDPC_TABLE_DATA_WIDTH)),
    3272 => std_logic_vector(to_unsigned(413, LDPC_TABLE_DATA_WIDTH)),
    3273 => std_logic_vector(to_unsigned(4455, LDPC_TABLE_DATA_WIDTH)),
    3274 => std_logic_vector(to_unsigned(2262, LDPC_TABLE_DATA_WIDTH)),
    3275 => std_logic_vector(to_unsigned(7915, LDPC_TABLE_DATA_WIDTH)),
    3276 => std_logic_vector(to_unsigned(12402, LDPC_TABLE_DATA_WIDTH)),
    3277 => std_logic_vector(to_unsigned(8579, LDPC_TABLE_DATA_WIDTH)),
    3278 => std_logic_vector(to_unsigned(7052, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3279 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    3280 => std_logic_vector(to_unsigned(3885, LDPC_TABLE_DATA_WIDTH)),
    3281 => std_logic_vector(to_unsigned(9126, LDPC_TABLE_DATA_WIDTH)),
    3282 => std_logic_vector(to_unsigned(5665, LDPC_TABLE_DATA_WIDTH)),
    3283 => std_logic_vector(to_unsigned(4505, LDPC_TABLE_DATA_WIDTH)),
    3284 => std_logic_vector(to_unsigned(2343, LDPC_TABLE_DATA_WIDTH)),
    3285 => std_logic_vector(to_unsigned(253, LDPC_TABLE_DATA_WIDTH)),
    3286 => std_logic_vector(to_unsigned(4707, LDPC_TABLE_DATA_WIDTH)),
    3287 => std_logic_vector(to_unsigned(3742, LDPC_TABLE_DATA_WIDTH)),
    3288 => std_logic_vector(to_unsigned(4166, LDPC_TABLE_DATA_WIDTH)),
    3289 => std_logic_vector(to_unsigned(1556, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3290 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    3291 => std_logic_vector(to_unsigned(1704, LDPC_TABLE_DATA_WIDTH)),
    3292 => std_logic_vector(to_unsigned(8936, LDPC_TABLE_DATA_WIDTH)),
    3293 => std_logic_vector(to_unsigned(6775, LDPC_TABLE_DATA_WIDTH)),
    3294 => std_logic_vector(to_unsigned(8639, LDPC_TABLE_DATA_WIDTH)),
    3295 => std_logic_vector(to_unsigned(8179, LDPC_TABLE_DATA_WIDTH)),
    3296 => std_logic_vector(to_unsigned(7954, LDPC_TABLE_DATA_WIDTH)),
    3297 => std_logic_vector(to_unsigned(8234, LDPC_TABLE_DATA_WIDTH)),
    3298 => std_logic_vector(to_unsigned(7850, LDPC_TABLE_DATA_WIDTH)),
    3299 => std_logic_vector(to_unsigned(8883, LDPC_TABLE_DATA_WIDTH)),
    3300 => std_logic_vector(to_unsigned(8713, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3301 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    3302 => std_logic_vector(to_unsigned(11716, LDPC_TABLE_DATA_WIDTH)),
    3303 => std_logic_vector(to_unsigned(4344, LDPC_TABLE_DATA_WIDTH)),
    3304 => std_logic_vector(to_unsigned(9087, LDPC_TABLE_DATA_WIDTH)),
    3305 => std_logic_vector(to_unsigned(11264, LDPC_TABLE_DATA_WIDTH)),
    3306 => std_logic_vector(to_unsigned(2274, LDPC_TABLE_DATA_WIDTH)),
    3307 => std_logic_vector(to_unsigned(8832, LDPC_TABLE_DATA_WIDTH)),
    3308 => std_logic_vector(to_unsigned(9147, LDPC_TABLE_DATA_WIDTH)),
    3309 => std_logic_vector(to_unsigned(11930, LDPC_TABLE_DATA_WIDTH)),
    3310 => std_logic_vector(to_unsigned(6054, LDPC_TABLE_DATA_WIDTH)),
    3311 => std_logic_vector(to_unsigned(5455, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3312 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3313 => std_logic_vector(to_unsigned(7323, LDPC_TABLE_DATA_WIDTH)),
    3314 => std_logic_vector(to_unsigned(3970, LDPC_TABLE_DATA_WIDTH)),
    3315 => std_logic_vector(to_unsigned(10329, LDPC_TABLE_DATA_WIDTH)),
    3316 => std_logic_vector(to_unsigned(2170, LDPC_TABLE_DATA_WIDTH)),
    3317 => std_logic_vector(to_unsigned(8262, LDPC_TABLE_DATA_WIDTH)),
    3318 => std_logic_vector(to_unsigned(3854, LDPC_TABLE_DATA_WIDTH)),
    3319 => std_logic_vector(to_unsigned(2087, LDPC_TABLE_DATA_WIDTH)),
    3320 => std_logic_vector(to_unsigned(12899, LDPC_TABLE_DATA_WIDTH)),
    3321 => std_logic_vector(to_unsigned(9497, LDPC_TABLE_DATA_WIDTH)),
    3322 => std_logic_vector(to_unsigned(11700, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3323 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3324 => std_logic_vector(to_unsigned(4418, LDPC_TABLE_DATA_WIDTH)),
    3325 => std_logic_vector(to_unsigned(1467, LDPC_TABLE_DATA_WIDTH)),
    3326 => std_logic_vector(to_unsigned(2490, LDPC_TABLE_DATA_WIDTH)),
    3327 => std_logic_vector(to_unsigned(5841, LDPC_TABLE_DATA_WIDTH)),
    3328 => std_logic_vector(to_unsigned(817, LDPC_TABLE_DATA_WIDTH)),
    3329 => std_logic_vector(to_unsigned(11453, LDPC_TABLE_DATA_WIDTH)),
    3330 => std_logic_vector(to_unsigned(533, LDPC_TABLE_DATA_WIDTH)),
    3331 => std_logic_vector(to_unsigned(11217, LDPC_TABLE_DATA_WIDTH)),
    3332 => std_logic_vector(to_unsigned(11962, LDPC_TABLE_DATA_WIDTH)),
    3333 => std_logic_vector(to_unsigned(5251, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3334 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3335 => std_logic_vector(to_unsigned(1541, LDPC_TABLE_DATA_WIDTH)),
    3336 => std_logic_vector(to_unsigned(4525, LDPC_TABLE_DATA_WIDTH)),
    3337 => std_logic_vector(to_unsigned(7976, LDPC_TABLE_DATA_WIDTH)),
    3338 => std_logic_vector(to_unsigned(3457, LDPC_TABLE_DATA_WIDTH)),
    3339 => std_logic_vector(to_unsigned(9536, LDPC_TABLE_DATA_WIDTH)),
    3340 => std_logic_vector(to_unsigned(7725, LDPC_TABLE_DATA_WIDTH)),
    3341 => std_logic_vector(to_unsigned(3788, LDPC_TABLE_DATA_WIDTH)),
    3342 => std_logic_vector(to_unsigned(2982, LDPC_TABLE_DATA_WIDTH)),
    3343 => std_logic_vector(to_unsigned(6307, LDPC_TABLE_DATA_WIDTH)),
    3344 => std_logic_vector(to_unsigned(5997, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3345 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3346 => std_logic_vector(to_unsigned(11484, LDPC_TABLE_DATA_WIDTH)),
    3347 => std_logic_vector(to_unsigned(2739, LDPC_TABLE_DATA_WIDTH)),
    3348 => std_logic_vector(to_unsigned(4023, LDPC_TABLE_DATA_WIDTH)),
    3349 => std_logic_vector(to_unsigned(12107, LDPC_TABLE_DATA_WIDTH)),
    3350 => std_logic_vector(to_unsigned(6516, LDPC_TABLE_DATA_WIDTH)),
    3351 => std_logic_vector(to_unsigned(551, LDPC_TABLE_DATA_WIDTH)),
    3352 => std_logic_vector(to_unsigned(2572, LDPC_TABLE_DATA_WIDTH)),
    3353 => std_logic_vector(to_unsigned(6628, LDPC_TABLE_DATA_WIDTH)),
    3354 => std_logic_vector(to_unsigned(8150, LDPC_TABLE_DATA_WIDTH)),
    3355 => std_logic_vector(to_unsigned(9852, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3356 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3357 => std_logic_vector(to_unsigned(6070, LDPC_TABLE_DATA_WIDTH)),
    3358 => std_logic_vector(to_unsigned(1761, LDPC_TABLE_DATA_WIDTH)),
    3359 => std_logic_vector(to_unsigned(4627, LDPC_TABLE_DATA_WIDTH)),
    3360 => std_logic_vector(to_unsigned(6534, LDPC_TABLE_DATA_WIDTH)),
    3361 => std_logic_vector(to_unsigned(7913, LDPC_TABLE_DATA_WIDTH)),
    3362 => std_logic_vector(to_unsigned(3730, LDPC_TABLE_DATA_WIDTH)),
    3363 => std_logic_vector(to_unsigned(11866, LDPC_TABLE_DATA_WIDTH)),
    3364 => std_logic_vector(to_unsigned(1813, LDPC_TABLE_DATA_WIDTH)),
    3365 => std_logic_vector(to_unsigned(12306, LDPC_TABLE_DATA_WIDTH)),
    3366 => std_logic_vector(to_unsigned(8249, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3367 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3368 => std_logic_vector(to_unsigned(12441, LDPC_TABLE_DATA_WIDTH)),
    3369 => std_logic_vector(to_unsigned(5489, LDPC_TABLE_DATA_WIDTH)),
    3370 => std_logic_vector(to_unsigned(8748, LDPC_TABLE_DATA_WIDTH)),
    3371 => std_logic_vector(to_unsigned(7837, LDPC_TABLE_DATA_WIDTH)),
    3372 => std_logic_vector(to_unsigned(7660, LDPC_TABLE_DATA_WIDTH)),
    3373 => std_logic_vector(to_unsigned(2102, LDPC_TABLE_DATA_WIDTH)),
    3374 => std_logic_vector(to_unsigned(11341, LDPC_TABLE_DATA_WIDTH)),
    3375 => std_logic_vector(to_unsigned(2936, LDPC_TABLE_DATA_WIDTH)),
    3376 => std_logic_vector(to_unsigned(6712, LDPC_TABLE_DATA_WIDTH)),
    3377 => std_logic_vector(to_unsigned(11977, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3378 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3379 => std_logic_vector(to_unsigned(10155, LDPC_TABLE_DATA_WIDTH)),
    3380 => std_logic_vector(to_unsigned(4210, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3381 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3382 => std_logic_vector(to_unsigned(1010, LDPC_TABLE_DATA_WIDTH)),
    3383 => std_logic_vector(to_unsigned(10483, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3384 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3385 => std_logic_vector(to_unsigned(8900, LDPC_TABLE_DATA_WIDTH)),
    3386 => std_logic_vector(to_unsigned(10250, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3387 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3388 => std_logic_vector(to_unsigned(10243, LDPC_TABLE_DATA_WIDTH)),
    3389 => std_logic_vector(to_unsigned(12278, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3390 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3391 => std_logic_vector(to_unsigned(7070, LDPC_TABLE_DATA_WIDTH)),
    3392 => std_logic_vector(to_unsigned(4397, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3393 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3394 => std_logic_vector(to_unsigned(12271, LDPC_TABLE_DATA_WIDTH)),
    3395 => std_logic_vector(to_unsigned(3887, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3396 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3397 => std_logic_vector(to_unsigned(11980, LDPC_TABLE_DATA_WIDTH)),
    3398 => std_logic_vector(to_unsigned(6836, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3399 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3400 => std_logic_vector(to_unsigned(9514, LDPC_TABLE_DATA_WIDTH)),
    3401 => std_logic_vector(to_unsigned(4356, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3402 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3403 => std_logic_vector(to_unsigned(7137, LDPC_TABLE_DATA_WIDTH)),
    3404 => std_logic_vector(to_unsigned(10281, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3405 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3406 => std_logic_vector(to_unsigned(11881, LDPC_TABLE_DATA_WIDTH)),
    3407 => std_logic_vector(to_unsigned(2526, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3408 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3409 => std_logic_vector(to_unsigned(1969, LDPC_TABLE_DATA_WIDTH)),
    3410 => std_logic_vector(to_unsigned(11477, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3411 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3412 => std_logic_vector(to_unsigned(3044, LDPC_TABLE_DATA_WIDTH)),
    3413 => std_logic_vector(to_unsigned(10921, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3414 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    3415 => std_logic_vector(to_unsigned(2236, LDPC_TABLE_DATA_WIDTH)),
    3416 => std_logic_vector(to_unsigned(8724, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3417 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    3418 => std_logic_vector(to_unsigned(9104, LDPC_TABLE_DATA_WIDTH)),
    3419 => std_logic_vector(to_unsigned(6340, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3420 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    3421 => std_logic_vector(to_unsigned(7342, LDPC_TABLE_DATA_WIDTH)),
    3422 => std_logic_vector(to_unsigned(8582, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3423 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    3424 => std_logic_vector(to_unsigned(11675, LDPC_TABLE_DATA_WIDTH)),
    3425 => std_logic_vector(to_unsigned(10405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3426 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    3427 => std_logic_vector(to_unsigned(6467, LDPC_TABLE_DATA_WIDTH)),
    3428 => std_logic_vector(to_unsigned(12775, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3429 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    3430 => std_logic_vector(to_unsigned(3186, LDPC_TABLE_DATA_WIDTH)),
    3431 => std_logic_vector(to_unsigned(12198, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3432 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3433 => std_logic_vector(to_unsigned(9621, LDPC_TABLE_DATA_WIDTH)),
    3434 => std_logic_vector(to_unsigned(11445, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3435 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    3436 => std_logic_vector(to_unsigned(7486, LDPC_TABLE_DATA_WIDTH)),
    3437 => std_logic_vector(to_unsigned(5611, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3438 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    3439 => std_logic_vector(to_unsigned(4319, LDPC_TABLE_DATA_WIDTH)),
    3440 => std_logic_vector(to_unsigned(4879, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3441 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    3442 => std_logic_vector(to_unsigned(2196, LDPC_TABLE_DATA_WIDTH)),
    3443 => std_logic_vector(to_unsigned(344, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3444 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    3445 => std_logic_vector(to_unsigned(7527, LDPC_TABLE_DATA_WIDTH)),
    3446 => std_logic_vector(to_unsigned(6650, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3447 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    3448 => std_logic_vector(to_unsigned(10693, LDPC_TABLE_DATA_WIDTH)),
    3449 => std_logic_vector(to_unsigned(2440, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3450 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    3451 => std_logic_vector(to_unsigned(6755, LDPC_TABLE_DATA_WIDTH)),
    3452 => std_logic_vector(to_unsigned(2706, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3453 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    3454 => std_logic_vector(to_unsigned(5144, LDPC_TABLE_DATA_WIDTH)),
    3455 => std_logic_vector(to_unsigned(5998, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3456 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    3457 => std_logic_vector(to_unsigned(11043, LDPC_TABLE_DATA_WIDTH)),
    3458 => std_logic_vector(to_unsigned(8033, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3459 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    3460 => std_logic_vector(to_unsigned(4846, LDPC_TABLE_DATA_WIDTH)),
    3461 => std_logic_vector(to_unsigned(4435, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3462 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    3463 => std_logic_vector(to_unsigned(4157, LDPC_TABLE_DATA_WIDTH)),
    3464 => std_logic_vector(to_unsigned(9228, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3465 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    3466 => std_logic_vector(to_unsigned(12270, LDPC_TABLE_DATA_WIDTH)),
    3467 => std_logic_vector(to_unsigned(6562, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3468 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3469 => std_logic_vector(to_unsigned(11954, LDPC_TABLE_DATA_WIDTH)),
    3470 => std_logic_vector(to_unsigned(7592, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3471 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3472 => std_logic_vector(to_unsigned(7420, LDPC_TABLE_DATA_WIDTH)),
    3473 => std_logic_vector(to_unsigned(2592, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3474 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3475 => std_logic_vector(to_unsigned(8810, LDPC_TABLE_DATA_WIDTH)),
    3476 => std_logic_vector(to_unsigned(9636, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3477 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3478 => std_logic_vector(to_unsigned(689, LDPC_TABLE_DATA_WIDTH)),
    3479 => std_logic_vector(to_unsigned(5430, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3480 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3481 => std_logic_vector(to_unsigned(920, LDPC_TABLE_DATA_WIDTH)),
    3482 => std_logic_vector(to_unsigned(1304, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3483 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3484 => std_logic_vector(to_unsigned(1253, LDPC_TABLE_DATA_WIDTH)),
    3485 => std_logic_vector(to_unsigned(11934, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3486 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3487 => std_logic_vector(to_unsigned(9559, LDPC_TABLE_DATA_WIDTH)),
    3488 => std_logic_vector(to_unsigned(6016, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3489 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3490 => std_logic_vector(to_unsigned(312, LDPC_TABLE_DATA_WIDTH)),
    3491 => std_logic_vector(to_unsigned(7589, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3492 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3493 => std_logic_vector(to_unsigned(4439, LDPC_TABLE_DATA_WIDTH)),
    3494 => std_logic_vector(to_unsigned(4197, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3495 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3496 => std_logic_vector(to_unsigned(4002, LDPC_TABLE_DATA_WIDTH)),
    3497 => std_logic_vector(to_unsigned(9555, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3498 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3499 => std_logic_vector(to_unsigned(12232, LDPC_TABLE_DATA_WIDTH)),
    3500 => std_logic_vector(to_unsigned(7779, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3501 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3502 => std_logic_vector(to_unsigned(1494, LDPC_TABLE_DATA_WIDTH)),
    3503 => std_logic_vector(to_unsigned(8782, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3504 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3505 => std_logic_vector(to_unsigned(10749, LDPC_TABLE_DATA_WIDTH)),
    3506 => std_logic_vector(to_unsigned(3969, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3507 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3508 => std_logic_vector(to_unsigned(4368, LDPC_TABLE_DATA_WIDTH)),
    3509 => std_logic_vector(to_unsigned(3479, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3510 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3511 => std_logic_vector(to_unsigned(6316, LDPC_TABLE_DATA_WIDTH)),
    3512 => std_logic_vector(to_unsigned(5342, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3513 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3514 => std_logic_vector(to_unsigned(2455, LDPC_TABLE_DATA_WIDTH)),
    3515 => std_logic_vector(to_unsigned(3493, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3516 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3517 => std_logic_vector(to_unsigned(12157, LDPC_TABLE_DATA_WIDTH)),
    3518 => std_logic_vector(to_unsigned(7405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3519 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3520 => std_logic_vector(to_unsigned(6598, LDPC_TABLE_DATA_WIDTH)),
    3521 => std_logic_vector(to_unsigned(11495, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3522 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    3523 => std_logic_vector(to_unsigned(11805, LDPC_TABLE_DATA_WIDTH)),
    3524 => std_logic_vector(to_unsigned(4455, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3525 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    3526 => std_logic_vector(to_unsigned(9625, LDPC_TABLE_DATA_WIDTH)),
    3527 => std_logic_vector(to_unsigned(2090, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3528 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    3529 => std_logic_vector(to_unsigned(4731, LDPC_TABLE_DATA_WIDTH)),
    3530 => std_logic_vector(to_unsigned(2321, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3531 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    3532 => std_logic_vector(to_unsigned(3578, LDPC_TABLE_DATA_WIDTH)),
    3533 => std_logic_vector(to_unsigned(2608, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3534 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    3535 => std_logic_vector(to_unsigned(8504, LDPC_TABLE_DATA_WIDTH)),
    3536 => std_logic_vector(to_unsigned(1849, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3537 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    3538 => std_logic_vector(to_unsigned(4027, LDPC_TABLE_DATA_WIDTH)),
    3539 => std_logic_vector(to_unsigned(1151, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3540 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3541 => std_logic_vector(to_unsigned(5647, LDPC_TABLE_DATA_WIDTH)),
    3542 => std_logic_vector(to_unsigned(4935, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3543 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    3544 => std_logic_vector(to_unsigned(4219, LDPC_TABLE_DATA_WIDTH)),
    3545 => std_logic_vector(to_unsigned(1870, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3546 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    3547 => std_logic_vector(to_unsigned(10968, LDPC_TABLE_DATA_WIDTH)),
    3548 => std_logic_vector(to_unsigned(8054, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3549 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    3550 => std_logic_vector(to_unsigned(6970, LDPC_TABLE_DATA_WIDTH)),
    3551 => std_logic_vector(to_unsigned(5447, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3552 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    3553 => std_logic_vector(to_unsigned(3217, LDPC_TABLE_DATA_WIDTH)),
    3554 => std_logic_vector(to_unsigned(5638, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3555 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    3556 => std_logic_vector(to_unsigned(8972, LDPC_TABLE_DATA_WIDTH)),
    3557 => std_logic_vector(to_unsigned(669, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3558 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    3559 => std_logic_vector(to_unsigned(5618, LDPC_TABLE_DATA_WIDTH)),
    3560 => std_logic_vector(to_unsigned(12472, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3561 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    3562 => std_logic_vector(to_unsigned(1457, LDPC_TABLE_DATA_WIDTH)),
    3563 => std_logic_vector(to_unsigned(1280, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3564 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    3565 => std_logic_vector(to_unsigned(8868, LDPC_TABLE_DATA_WIDTH)),
    3566 => std_logic_vector(to_unsigned(3883, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3567 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    3568 => std_logic_vector(to_unsigned(8866, LDPC_TABLE_DATA_WIDTH)),
    3569 => std_logic_vector(to_unsigned(1224, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3570 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    3571 => std_logic_vector(to_unsigned(8371, LDPC_TABLE_DATA_WIDTH)),
    3572 => std_logic_vector(to_unsigned(5972, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3573 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    3574 => std_logic_vector(to_unsigned(266, LDPC_TABLE_DATA_WIDTH)),
    3575 => std_logic_vector(to_unsigned(4405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3576 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3577 => std_logic_vector(to_unsigned(3706, LDPC_TABLE_DATA_WIDTH)),
    3578 => std_logic_vector(to_unsigned(3244, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3579 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3580 => std_logic_vector(to_unsigned(6039, LDPC_TABLE_DATA_WIDTH)),
    3581 => std_logic_vector(to_unsigned(5844, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3582 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3583 => std_logic_vector(to_unsigned(7200, LDPC_TABLE_DATA_WIDTH)),
    3584 => std_logic_vector(to_unsigned(3283, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3585 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3586 => std_logic_vector(to_unsigned(1502, LDPC_TABLE_DATA_WIDTH)),
    3587 => std_logic_vector(to_unsigned(11282, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3588 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3589 => std_logic_vector(to_unsigned(12318, LDPC_TABLE_DATA_WIDTH)),
    3590 => std_logic_vector(to_unsigned(2202, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3591 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3592 => std_logic_vector(to_unsigned(4523, LDPC_TABLE_DATA_WIDTH)),
    3593 => std_logic_vector(to_unsigned(965, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3594 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3595 => std_logic_vector(to_unsigned(9587, LDPC_TABLE_DATA_WIDTH)),
    3596 => std_logic_vector(to_unsigned(7011, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3597 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3598 => std_logic_vector(to_unsigned(2552, LDPC_TABLE_DATA_WIDTH)),
    3599 => std_logic_vector(to_unsigned(2051, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3600 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3601 => std_logic_vector(to_unsigned(12045, LDPC_TABLE_DATA_WIDTH)),
    3602 => std_logic_vector(to_unsigned(10306, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3603 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3604 => std_logic_vector(to_unsigned(11070, LDPC_TABLE_DATA_WIDTH)),
    3605 => std_logic_vector(to_unsigned(5104, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3606 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3607 => std_logic_vector(to_unsigned(6627, LDPC_TABLE_DATA_WIDTH)),
    3608 => std_logic_vector(to_unsigned(6906, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3609 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3610 => std_logic_vector(to_unsigned(9889, LDPC_TABLE_DATA_WIDTH)),
    3611 => std_logic_vector(to_unsigned(2121, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3612 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3613 => std_logic_vector(to_unsigned(829, LDPC_TABLE_DATA_WIDTH)),
    3614 => std_logic_vector(to_unsigned(9701, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3615 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3616 => std_logic_vector(to_unsigned(2201, LDPC_TABLE_DATA_WIDTH)),
    3617 => std_logic_vector(to_unsigned(1819, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3618 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3619 => std_logic_vector(to_unsigned(6689, LDPC_TABLE_DATA_WIDTH)),
    3620 => std_logic_vector(to_unsigned(12925, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3621 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3622 => std_logic_vector(to_unsigned(2139, LDPC_TABLE_DATA_WIDTH)),
    3623 => std_logic_vector(to_unsigned(8757, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3624 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3625 => std_logic_vector(to_unsigned(12004, LDPC_TABLE_DATA_WIDTH)),
    3626 => std_logic_vector(to_unsigned(5948, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3627 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3628 => std_logic_vector(to_unsigned(8704, LDPC_TABLE_DATA_WIDTH)),
    3629 => std_logic_vector(to_unsigned(3191, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3630 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    3631 => std_logic_vector(to_unsigned(8171, LDPC_TABLE_DATA_WIDTH)),
    3632 => std_logic_vector(to_unsigned(10933, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3633 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    3634 => std_logic_vector(to_unsigned(6297, LDPC_TABLE_DATA_WIDTH)),
    3635 => std_logic_vector(to_unsigned(7116, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3636 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    3637 => std_logic_vector(to_unsigned(616, LDPC_TABLE_DATA_WIDTH)),
    3638 => std_logic_vector(to_unsigned(7146, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3639 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    3640 => std_logic_vector(to_unsigned(5142, LDPC_TABLE_DATA_WIDTH)),
    3641 => std_logic_vector(to_unsigned(9761, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3642 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    3643 => std_logic_vector(to_unsigned(10377, LDPC_TABLE_DATA_WIDTH)),
    3644 => std_logic_vector(to_unsigned(8138, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3645 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    3646 => std_logic_vector(to_unsigned(7616, LDPC_TABLE_DATA_WIDTH)),
    3647 => std_logic_vector(to_unsigned(5811, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3648 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3649 => std_logic_vector(to_unsigned(7285, LDPC_TABLE_DATA_WIDTH)),
    3650 => std_logic_vector(to_unsigned(9863, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3651 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    3652 => std_logic_vector(to_unsigned(7764, LDPC_TABLE_DATA_WIDTH)),
    3653 => std_logic_vector(to_unsigned(10867, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3654 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    3655 => std_logic_vector(to_unsigned(12343, LDPC_TABLE_DATA_WIDTH)),
    3656 => std_logic_vector(to_unsigned(9019, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3657 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    3658 => std_logic_vector(to_unsigned(4414, LDPC_TABLE_DATA_WIDTH)),
    3659 => std_logic_vector(to_unsigned(8331, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3660 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    3661 => std_logic_vector(to_unsigned(3464, LDPC_TABLE_DATA_WIDTH)),
    3662 => std_logic_vector(to_unsigned(642, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3663 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    3664 => std_logic_vector(to_unsigned(6960, LDPC_TABLE_DATA_WIDTH)),
    3665 => std_logic_vector(to_unsigned(2039, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3666 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    3667 => std_logic_vector(to_unsigned(786, LDPC_TABLE_DATA_WIDTH)),
    3668 => std_logic_vector(to_unsigned(3021, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3669 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    3670 => std_logic_vector(to_unsigned(710, LDPC_TABLE_DATA_WIDTH)),
    3671 => std_logic_vector(to_unsigned(2086, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3672 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    3673 => std_logic_vector(to_unsigned(7423, LDPC_TABLE_DATA_WIDTH)),
    3674 => std_logic_vector(to_unsigned(5601, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3675 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    3676 => std_logic_vector(to_unsigned(8120, LDPC_TABLE_DATA_WIDTH)),
    3677 => std_logic_vector(to_unsigned(4885, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3678 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    3679 => std_logic_vector(to_unsigned(12385, LDPC_TABLE_DATA_WIDTH)),
    3680 => std_logic_vector(to_unsigned(11990, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3681 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    3682 => std_logic_vector(to_unsigned(9739, LDPC_TABLE_DATA_WIDTH)),
    3683 => std_logic_vector(to_unsigned(10034, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3684 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3685 => std_logic_vector(to_unsigned(424, LDPC_TABLE_DATA_WIDTH)),
    3686 => std_logic_vector(to_unsigned(10162, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3687 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3688 => std_logic_vector(to_unsigned(1347, LDPC_TABLE_DATA_WIDTH)),
    3689 => std_logic_vector(to_unsigned(7597, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3690 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3691 => std_logic_vector(to_unsigned(1450, LDPC_TABLE_DATA_WIDTH)),
    3692 => std_logic_vector(to_unsigned(112, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3693 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3694 => std_logic_vector(to_unsigned(7965, LDPC_TABLE_DATA_WIDTH)),
    3695 => std_logic_vector(to_unsigned(8478, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3696 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3697 => std_logic_vector(to_unsigned(8945, LDPC_TABLE_DATA_WIDTH)),
    3698 => std_logic_vector(to_unsigned(7397, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3699 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3700 => std_logic_vector(to_unsigned(6590, LDPC_TABLE_DATA_WIDTH)),
    3701 => std_logic_vector(to_unsigned(8316, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3702 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3703 => std_logic_vector(to_unsigned(6838, LDPC_TABLE_DATA_WIDTH)),
    3704 => std_logic_vector(to_unsigned(9011, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3705 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3706 => std_logic_vector(to_unsigned(6174, LDPC_TABLE_DATA_WIDTH)),
    3707 => std_logic_vector(to_unsigned(9410, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3708 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3709 => std_logic_vector(to_unsigned(255, LDPC_TABLE_DATA_WIDTH)),
    3710 => std_logic_vector(to_unsigned(113, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3711 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3712 => std_logic_vector(to_unsigned(6197, LDPC_TABLE_DATA_WIDTH)),
    3713 => std_logic_vector(to_unsigned(5835, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3714 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3715 => std_logic_vector(to_unsigned(12902, LDPC_TABLE_DATA_WIDTH)),
    3716 => std_logic_vector(to_unsigned(3844, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3717 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3718 => std_logic_vector(to_unsigned(4377, LDPC_TABLE_DATA_WIDTH)),
    3719 => std_logic_vector(to_unsigned(3505, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3720 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3721 => std_logic_vector(to_unsigned(5478, LDPC_TABLE_DATA_WIDTH)),
    3722 => std_logic_vector(to_unsigned(8672, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3723 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3724 => std_logic_vector(to_unsigned(4453, LDPC_TABLE_DATA_WIDTH)),
    3725 => std_logic_vector(to_unsigned(2132, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3726 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3727 => std_logic_vector(to_unsigned(9724, LDPC_TABLE_DATA_WIDTH)),
    3728 => std_logic_vector(to_unsigned(1380, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3729 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3730 => std_logic_vector(to_unsigned(12131, LDPC_TABLE_DATA_WIDTH)),
    3731 => std_logic_vector(to_unsigned(11526, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3732 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3733 => std_logic_vector(to_unsigned(12323, LDPC_TABLE_DATA_WIDTH)),
    3734 => std_logic_vector(to_unsigned(9511, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3735 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3736 => std_logic_vector(to_unsigned(8231, LDPC_TABLE_DATA_WIDTH)),
    3737 => std_logic_vector(to_unsigned(1752, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3738 => std_logic_vector(to_unsigned(30, LDPC_TABLE_DATA_WIDTH)),
    3739 => std_logic_vector(to_unsigned(497, LDPC_TABLE_DATA_WIDTH)),
    3740 => std_logic_vector(to_unsigned(9022, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3741 => std_logic_vector(to_unsigned(31, LDPC_TABLE_DATA_WIDTH)),
    3742 => std_logic_vector(to_unsigned(9288, LDPC_TABLE_DATA_WIDTH)),
    3743 => std_logic_vector(to_unsigned(3080, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3744 => std_logic_vector(to_unsigned(32, LDPC_TABLE_DATA_WIDTH)),
    3745 => std_logic_vector(to_unsigned(2481, LDPC_TABLE_DATA_WIDTH)),
    3746 => std_logic_vector(to_unsigned(7515, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3747 => std_logic_vector(to_unsigned(33, LDPC_TABLE_DATA_WIDTH)),
    3748 => std_logic_vector(to_unsigned(2696, LDPC_TABLE_DATA_WIDTH)),
    3749 => std_logic_vector(to_unsigned(268, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3750 => std_logic_vector(to_unsigned(34, LDPC_TABLE_DATA_WIDTH)),
    3751 => std_logic_vector(to_unsigned(4023, LDPC_TABLE_DATA_WIDTH)),
    3752 => std_logic_vector(to_unsigned(12341, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3753 => std_logic_vector(to_unsigned(35, LDPC_TABLE_DATA_WIDTH)),
    3754 => std_logic_vector(to_unsigned(7108, LDPC_TABLE_DATA_WIDTH)),
    3755 => std_logic_vector(to_unsigned(5553, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C5_6
    3756 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3757 => std_logic_vector(to_unsigned(4362, LDPC_TABLE_DATA_WIDTH)),
    3758 => std_logic_vector(to_unsigned(416, LDPC_TABLE_DATA_WIDTH)),
    3759 => std_logic_vector(to_unsigned(8909, LDPC_TABLE_DATA_WIDTH)),
    3760 => std_logic_vector(to_unsigned(4156, LDPC_TABLE_DATA_WIDTH)),
    3761 => std_logic_vector(to_unsigned(3216, LDPC_TABLE_DATA_WIDTH)),
    3762 => std_logic_vector(to_unsigned(3112, LDPC_TABLE_DATA_WIDTH)),
    3763 => std_logic_vector(to_unsigned(2560, LDPC_TABLE_DATA_WIDTH)),
    3764 => std_logic_vector(to_unsigned(2912, LDPC_TABLE_DATA_WIDTH)),
    3765 => std_logic_vector(to_unsigned(6405, LDPC_TABLE_DATA_WIDTH)),
    3766 => std_logic_vector(to_unsigned(8593, LDPC_TABLE_DATA_WIDTH)),
    3767 => std_logic_vector(to_unsigned(4969, LDPC_TABLE_DATA_WIDTH)),
    3768 => std_logic_vector(to_unsigned(6723, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3769 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    3770 => std_logic_vector(to_unsigned(2479, LDPC_TABLE_DATA_WIDTH)),
    3771 => std_logic_vector(to_unsigned(1786, LDPC_TABLE_DATA_WIDTH)),
    3772 => std_logic_vector(to_unsigned(8978, LDPC_TABLE_DATA_WIDTH)),
    3773 => std_logic_vector(to_unsigned(3011, LDPC_TABLE_DATA_WIDTH)),
    3774 => std_logic_vector(to_unsigned(4339, LDPC_TABLE_DATA_WIDTH)),
    3775 => std_logic_vector(to_unsigned(9313, LDPC_TABLE_DATA_WIDTH)),
    3776 => std_logic_vector(to_unsigned(6397, LDPC_TABLE_DATA_WIDTH)),
    3777 => std_logic_vector(to_unsigned(2957, LDPC_TABLE_DATA_WIDTH)),
    3778 => std_logic_vector(to_unsigned(7288, LDPC_TABLE_DATA_WIDTH)),
    3779 => std_logic_vector(to_unsigned(5484, LDPC_TABLE_DATA_WIDTH)),
    3780 => std_logic_vector(to_unsigned(6031, LDPC_TABLE_DATA_WIDTH)),
    3781 => std_logic_vector(to_unsigned(10217, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3782 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    3783 => std_logic_vector(to_unsigned(10175, LDPC_TABLE_DATA_WIDTH)),
    3784 => std_logic_vector(to_unsigned(9009, LDPC_TABLE_DATA_WIDTH)),
    3785 => std_logic_vector(to_unsigned(9889, LDPC_TABLE_DATA_WIDTH)),
    3786 => std_logic_vector(to_unsigned(3091, LDPC_TABLE_DATA_WIDTH)),
    3787 => std_logic_vector(to_unsigned(4985, LDPC_TABLE_DATA_WIDTH)),
    3788 => std_logic_vector(to_unsigned(7267, LDPC_TABLE_DATA_WIDTH)),
    3789 => std_logic_vector(to_unsigned(4092, LDPC_TABLE_DATA_WIDTH)),
    3790 => std_logic_vector(to_unsigned(8874, LDPC_TABLE_DATA_WIDTH)),
    3791 => std_logic_vector(to_unsigned(5671, LDPC_TABLE_DATA_WIDTH)),
    3792 => std_logic_vector(to_unsigned(2777, LDPC_TABLE_DATA_WIDTH)),
    3793 => std_logic_vector(to_unsigned(2189, LDPC_TABLE_DATA_WIDTH)),
    3794 => std_logic_vector(to_unsigned(8716, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3795 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    3796 => std_logic_vector(to_unsigned(9052, LDPC_TABLE_DATA_WIDTH)),
    3797 => std_logic_vector(to_unsigned(4795, LDPC_TABLE_DATA_WIDTH)),
    3798 => std_logic_vector(to_unsigned(3924, LDPC_TABLE_DATA_WIDTH)),
    3799 => std_logic_vector(to_unsigned(3370, LDPC_TABLE_DATA_WIDTH)),
    3800 => std_logic_vector(to_unsigned(10058, LDPC_TABLE_DATA_WIDTH)),
    3801 => std_logic_vector(to_unsigned(1128, LDPC_TABLE_DATA_WIDTH)),
    3802 => std_logic_vector(to_unsigned(9996, LDPC_TABLE_DATA_WIDTH)),
    3803 => std_logic_vector(to_unsigned(10165, LDPC_TABLE_DATA_WIDTH)),
    3804 => std_logic_vector(to_unsigned(9360, LDPC_TABLE_DATA_WIDTH)),
    3805 => std_logic_vector(to_unsigned(4297, LDPC_TABLE_DATA_WIDTH)),
    3806 => std_logic_vector(to_unsigned(434, LDPC_TABLE_DATA_WIDTH)),
    3807 => std_logic_vector(to_unsigned(5138, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3808 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    3809 => std_logic_vector(to_unsigned(2379, LDPC_TABLE_DATA_WIDTH)),
    3810 => std_logic_vector(to_unsigned(7834, LDPC_TABLE_DATA_WIDTH)),
    3811 => std_logic_vector(to_unsigned(4835, LDPC_TABLE_DATA_WIDTH)),
    3812 => std_logic_vector(to_unsigned(2327, LDPC_TABLE_DATA_WIDTH)),
    3813 => std_logic_vector(to_unsigned(9843, LDPC_TABLE_DATA_WIDTH)),
    3814 => std_logic_vector(to_unsigned(804, LDPC_TABLE_DATA_WIDTH)),
    3815 => std_logic_vector(to_unsigned(329, LDPC_TABLE_DATA_WIDTH)),
    3816 => std_logic_vector(to_unsigned(8353, LDPC_TABLE_DATA_WIDTH)),
    3817 => std_logic_vector(to_unsigned(7167, LDPC_TABLE_DATA_WIDTH)),
    3818 => std_logic_vector(to_unsigned(3070, LDPC_TABLE_DATA_WIDTH)),
    3819 => std_logic_vector(to_unsigned(1528, LDPC_TABLE_DATA_WIDTH)),
    3820 => std_logic_vector(to_unsigned(7311, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3821 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    3822 => std_logic_vector(to_unsigned(3435, LDPC_TABLE_DATA_WIDTH)),
    3823 => std_logic_vector(to_unsigned(7871, LDPC_TABLE_DATA_WIDTH)),
    3824 => std_logic_vector(to_unsigned(348, LDPC_TABLE_DATA_WIDTH)),
    3825 => std_logic_vector(to_unsigned(3693, LDPC_TABLE_DATA_WIDTH)),
    3826 => std_logic_vector(to_unsigned(1876, LDPC_TABLE_DATA_WIDTH)),
    3827 => std_logic_vector(to_unsigned(6585, LDPC_TABLE_DATA_WIDTH)),
    3828 => std_logic_vector(to_unsigned(10340, LDPC_TABLE_DATA_WIDTH)),
    3829 => std_logic_vector(to_unsigned(7144, LDPC_TABLE_DATA_WIDTH)),
    3830 => std_logic_vector(to_unsigned(5870, LDPC_TABLE_DATA_WIDTH)),
    3831 => std_logic_vector(to_unsigned(2084, LDPC_TABLE_DATA_WIDTH)),
    3832 => std_logic_vector(to_unsigned(4052, LDPC_TABLE_DATA_WIDTH)),
    3833 => std_logic_vector(to_unsigned(2780, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3834 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    3835 => std_logic_vector(to_unsigned(3917, LDPC_TABLE_DATA_WIDTH)),
    3836 => std_logic_vector(to_unsigned(3111, LDPC_TABLE_DATA_WIDTH)),
    3837 => std_logic_vector(to_unsigned(3476, LDPC_TABLE_DATA_WIDTH)),
    3838 => std_logic_vector(to_unsigned(1304, LDPC_TABLE_DATA_WIDTH)),
    3839 => std_logic_vector(to_unsigned(10331, LDPC_TABLE_DATA_WIDTH)),
    3840 => std_logic_vector(to_unsigned(5939, LDPC_TABLE_DATA_WIDTH)),
    3841 => std_logic_vector(to_unsigned(5199, LDPC_TABLE_DATA_WIDTH)),
    3842 => std_logic_vector(to_unsigned(1611, LDPC_TABLE_DATA_WIDTH)),
    3843 => std_logic_vector(to_unsigned(1991, LDPC_TABLE_DATA_WIDTH)),
    3844 => std_logic_vector(to_unsigned(699, LDPC_TABLE_DATA_WIDTH)),
    3845 => std_logic_vector(to_unsigned(8316, LDPC_TABLE_DATA_WIDTH)),
    3846 => std_logic_vector(to_unsigned(9960, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3847 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    3848 => std_logic_vector(to_unsigned(6883, LDPC_TABLE_DATA_WIDTH)),
    3849 => std_logic_vector(to_unsigned(3237, LDPC_TABLE_DATA_WIDTH)),
    3850 => std_logic_vector(to_unsigned(1717, LDPC_TABLE_DATA_WIDTH)),
    3851 => std_logic_vector(to_unsigned(10752, LDPC_TABLE_DATA_WIDTH)),
    3852 => std_logic_vector(to_unsigned(7891, LDPC_TABLE_DATA_WIDTH)),
    3853 => std_logic_vector(to_unsigned(9764, LDPC_TABLE_DATA_WIDTH)),
    3854 => std_logic_vector(to_unsigned(4745, LDPC_TABLE_DATA_WIDTH)),
    3855 => std_logic_vector(to_unsigned(3888, LDPC_TABLE_DATA_WIDTH)),
    3856 => std_logic_vector(to_unsigned(10009, LDPC_TABLE_DATA_WIDTH)),
    3857 => std_logic_vector(to_unsigned(4176, LDPC_TABLE_DATA_WIDTH)),
    3858 => std_logic_vector(to_unsigned(4614, LDPC_TABLE_DATA_WIDTH)),
    3859 => std_logic_vector(to_unsigned(1567, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3860 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    3861 => std_logic_vector(to_unsigned(10587, LDPC_TABLE_DATA_WIDTH)),
    3862 => std_logic_vector(to_unsigned(2195, LDPC_TABLE_DATA_WIDTH)),
    3863 => std_logic_vector(to_unsigned(1689, LDPC_TABLE_DATA_WIDTH)),
    3864 => std_logic_vector(to_unsigned(2968, LDPC_TABLE_DATA_WIDTH)),
    3865 => std_logic_vector(to_unsigned(5420, LDPC_TABLE_DATA_WIDTH)),
    3866 => std_logic_vector(to_unsigned(2580, LDPC_TABLE_DATA_WIDTH)),
    3867 => std_logic_vector(to_unsigned(2883, LDPC_TABLE_DATA_WIDTH)),
    3868 => std_logic_vector(to_unsigned(6496, LDPC_TABLE_DATA_WIDTH)),
    3869 => std_logic_vector(to_unsigned(111, LDPC_TABLE_DATA_WIDTH)),
    3870 => std_logic_vector(to_unsigned(6023, LDPC_TABLE_DATA_WIDTH)),
    3871 => std_logic_vector(to_unsigned(1024, LDPC_TABLE_DATA_WIDTH)),
    3872 => std_logic_vector(to_unsigned(4449, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3873 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    3874 => std_logic_vector(to_unsigned(3786, LDPC_TABLE_DATA_WIDTH)),
    3875 => std_logic_vector(to_unsigned(8593, LDPC_TABLE_DATA_WIDTH)),
    3876 => std_logic_vector(to_unsigned(2074, LDPC_TABLE_DATA_WIDTH)),
    3877 => std_logic_vector(to_unsigned(3321, LDPC_TABLE_DATA_WIDTH)),
    3878 => std_logic_vector(to_unsigned(5057, LDPC_TABLE_DATA_WIDTH)),
    3879 => std_logic_vector(to_unsigned(1450, LDPC_TABLE_DATA_WIDTH)),
    3880 => std_logic_vector(to_unsigned(3840, LDPC_TABLE_DATA_WIDTH)),
    3881 => std_logic_vector(to_unsigned(5444, LDPC_TABLE_DATA_WIDTH)),
    3882 => std_logic_vector(to_unsigned(6572, LDPC_TABLE_DATA_WIDTH)),
    3883 => std_logic_vector(to_unsigned(3094, LDPC_TABLE_DATA_WIDTH)),
    3884 => std_logic_vector(to_unsigned(9892, LDPC_TABLE_DATA_WIDTH)),
    3885 => std_logic_vector(to_unsigned(1512, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3886 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    3887 => std_logic_vector(to_unsigned(8548, LDPC_TABLE_DATA_WIDTH)),
    3888 => std_logic_vector(to_unsigned(1848, LDPC_TABLE_DATA_WIDTH)),
    3889 => std_logic_vector(to_unsigned(10372, LDPC_TABLE_DATA_WIDTH)),
    3890 => std_logic_vector(to_unsigned(4585, LDPC_TABLE_DATA_WIDTH)),
    3891 => std_logic_vector(to_unsigned(7313, LDPC_TABLE_DATA_WIDTH)),
    3892 => std_logic_vector(to_unsigned(6536, LDPC_TABLE_DATA_WIDTH)),
    3893 => std_logic_vector(to_unsigned(6379, LDPC_TABLE_DATA_WIDTH)),
    3894 => std_logic_vector(to_unsigned(1766, LDPC_TABLE_DATA_WIDTH)),
    3895 => std_logic_vector(to_unsigned(9462, LDPC_TABLE_DATA_WIDTH)),
    3896 => std_logic_vector(to_unsigned(2456, LDPC_TABLE_DATA_WIDTH)),
    3897 => std_logic_vector(to_unsigned(5606, LDPC_TABLE_DATA_WIDTH)),
    3898 => std_logic_vector(to_unsigned(9975, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3899 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    3900 => std_logic_vector(to_unsigned(8204, LDPC_TABLE_DATA_WIDTH)),
    3901 => std_logic_vector(to_unsigned(10593, LDPC_TABLE_DATA_WIDTH)),
    3902 => std_logic_vector(to_unsigned(7935, LDPC_TABLE_DATA_WIDTH)),
    3903 => std_logic_vector(to_unsigned(3636, LDPC_TABLE_DATA_WIDTH)),
    3904 => std_logic_vector(to_unsigned(3882, LDPC_TABLE_DATA_WIDTH)),
    3905 => std_logic_vector(to_unsigned(394, LDPC_TABLE_DATA_WIDTH)),
    3906 => std_logic_vector(to_unsigned(5968, LDPC_TABLE_DATA_WIDTH)),
    3907 => std_logic_vector(to_unsigned(8561, LDPC_TABLE_DATA_WIDTH)),
    3908 => std_logic_vector(to_unsigned(2395, LDPC_TABLE_DATA_WIDTH)),
    3909 => std_logic_vector(to_unsigned(7289, LDPC_TABLE_DATA_WIDTH)),
    3910 => std_logic_vector(to_unsigned(9267, LDPC_TABLE_DATA_WIDTH)),
    3911 => std_logic_vector(to_unsigned(9978, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3912 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    3913 => std_logic_vector(to_unsigned(7795, LDPC_TABLE_DATA_WIDTH)),
    3914 => std_logic_vector(to_unsigned(74, LDPC_TABLE_DATA_WIDTH)),
    3915 => std_logic_vector(to_unsigned(1633, LDPC_TABLE_DATA_WIDTH)),
    3916 => std_logic_vector(to_unsigned(9542, LDPC_TABLE_DATA_WIDTH)),
    3917 => std_logic_vector(to_unsigned(6867, LDPC_TABLE_DATA_WIDTH)),
    3918 => std_logic_vector(to_unsigned(7352, LDPC_TABLE_DATA_WIDTH)),
    3919 => std_logic_vector(to_unsigned(6417, LDPC_TABLE_DATA_WIDTH)),
    3920 => std_logic_vector(to_unsigned(7568, LDPC_TABLE_DATA_WIDTH)),
    3921 => std_logic_vector(to_unsigned(10623, LDPC_TABLE_DATA_WIDTH)),
    3922 => std_logic_vector(to_unsigned(725, LDPC_TABLE_DATA_WIDTH)),
    3923 => std_logic_vector(to_unsigned(2531, LDPC_TABLE_DATA_WIDTH)),
    3924 => std_logic_vector(to_unsigned(9115, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3925 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    3926 => std_logic_vector(to_unsigned(7151, LDPC_TABLE_DATA_WIDTH)),
    3927 => std_logic_vector(to_unsigned(2482, LDPC_TABLE_DATA_WIDTH)),
    3928 => std_logic_vector(to_unsigned(4260, LDPC_TABLE_DATA_WIDTH)),
    3929 => std_logic_vector(to_unsigned(5003, LDPC_TABLE_DATA_WIDTH)),
    3930 => std_logic_vector(to_unsigned(10105, LDPC_TABLE_DATA_WIDTH)),
    3931 => std_logic_vector(to_unsigned(7419, LDPC_TABLE_DATA_WIDTH)),
    3932 => std_logic_vector(to_unsigned(9203, LDPC_TABLE_DATA_WIDTH)),
    3933 => std_logic_vector(to_unsigned(6691, LDPC_TABLE_DATA_WIDTH)),
    3934 => std_logic_vector(to_unsigned(8798, LDPC_TABLE_DATA_WIDTH)),
    3935 => std_logic_vector(to_unsigned(2092, LDPC_TABLE_DATA_WIDTH)),
    3936 => std_logic_vector(to_unsigned(8263, LDPC_TABLE_DATA_WIDTH)),
    3937 => std_logic_vector(to_unsigned(3755, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3938 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    3939 => std_logic_vector(to_unsigned(3600, LDPC_TABLE_DATA_WIDTH)),
    3940 => std_logic_vector(to_unsigned(570, LDPC_TABLE_DATA_WIDTH)),
    3941 => std_logic_vector(to_unsigned(4527, LDPC_TABLE_DATA_WIDTH)),
    3942 => std_logic_vector(to_unsigned(200, LDPC_TABLE_DATA_WIDTH)),
    3943 => std_logic_vector(to_unsigned(9718, LDPC_TABLE_DATA_WIDTH)),
    3944 => std_logic_vector(to_unsigned(6771, LDPC_TABLE_DATA_WIDTH)),
    3945 => std_logic_vector(to_unsigned(1995, LDPC_TABLE_DATA_WIDTH)),
    3946 => std_logic_vector(to_unsigned(8902, LDPC_TABLE_DATA_WIDTH)),
    3947 => std_logic_vector(to_unsigned(5446, LDPC_TABLE_DATA_WIDTH)),
    3948 => std_logic_vector(to_unsigned(768, LDPC_TABLE_DATA_WIDTH)),
    3949 => std_logic_vector(to_unsigned(1103, LDPC_TABLE_DATA_WIDTH)),
    3950 => std_logic_vector(to_unsigned(6520, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3951 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    3952 => std_logic_vector(to_unsigned(6304, LDPC_TABLE_DATA_WIDTH)),
    3953 => std_logic_vector(to_unsigned(7621, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3954 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    3955 => std_logic_vector(to_unsigned(6498, LDPC_TABLE_DATA_WIDTH)),
    3956 => std_logic_vector(to_unsigned(9209, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3957 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    3958 => std_logic_vector(to_unsigned(7293, LDPC_TABLE_DATA_WIDTH)),
    3959 => std_logic_vector(to_unsigned(6786, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3960 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    3961 => std_logic_vector(to_unsigned(5950, LDPC_TABLE_DATA_WIDTH)),
    3962 => std_logic_vector(to_unsigned(1708, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3963 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    3964 => std_logic_vector(to_unsigned(8521, LDPC_TABLE_DATA_WIDTH)),
    3965 => std_logic_vector(to_unsigned(1793, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3966 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    3967 => std_logic_vector(to_unsigned(6174, LDPC_TABLE_DATA_WIDTH)),
    3968 => std_logic_vector(to_unsigned(7854, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3969 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    3970 => std_logic_vector(to_unsigned(9773, LDPC_TABLE_DATA_WIDTH)),
    3971 => std_logic_vector(to_unsigned(1190, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3972 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    3973 => std_logic_vector(to_unsigned(9517, LDPC_TABLE_DATA_WIDTH)),
    3974 => std_logic_vector(to_unsigned(10268, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3975 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    3976 => std_logic_vector(to_unsigned(2181, LDPC_TABLE_DATA_WIDTH)),
    3977 => std_logic_vector(to_unsigned(9349, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3978 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    3979 => std_logic_vector(to_unsigned(1949, LDPC_TABLE_DATA_WIDTH)),
    3980 => std_logic_vector(to_unsigned(5560, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3981 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    3982 => std_logic_vector(to_unsigned(1556, LDPC_TABLE_DATA_WIDTH)),
    3983 => std_logic_vector(to_unsigned(555, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3984 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    3985 => std_logic_vector(to_unsigned(8600, LDPC_TABLE_DATA_WIDTH)),
    3986 => std_logic_vector(to_unsigned(3827, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3987 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    3988 => std_logic_vector(to_unsigned(5072, LDPC_TABLE_DATA_WIDTH)),
    3989 => std_logic_vector(to_unsigned(1057, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3990 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    3991 => std_logic_vector(to_unsigned(7928, LDPC_TABLE_DATA_WIDTH)),
    3992 => std_logic_vector(to_unsigned(3542, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3993 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    3994 => std_logic_vector(to_unsigned(3226, LDPC_TABLE_DATA_WIDTH)),
    3995 => std_logic_vector(to_unsigned(3762, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3996 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    3997 => std_logic_vector(to_unsigned(7045, LDPC_TABLE_DATA_WIDTH)),
    3998 => std_logic_vector(to_unsigned(2420, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    3999 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4000 => std_logic_vector(to_unsigned(9645, LDPC_TABLE_DATA_WIDTH)),
    4001 => std_logic_vector(to_unsigned(2641, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4002 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4003 => std_logic_vector(to_unsigned(2774, LDPC_TABLE_DATA_WIDTH)),
    4004 => std_logic_vector(to_unsigned(2452, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4005 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4006 => std_logic_vector(to_unsigned(5331, LDPC_TABLE_DATA_WIDTH)),
    4007 => std_logic_vector(to_unsigned(2031, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4008 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4009 => std_logic_vector(to_unsigned(9400, LDPC_TABLE_DATA_WIDTH)),
    4010 => std_logic_vector(to_unsigned(7503, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4011 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4012 => std_logic_vector(to_unsigned(1850, LDPC_TABLE_DATA_WIDTH)),
    4013 => std_logic_vector(to_unsigned(2338, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4014 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4015 => std_logic_vector(to_unsigned(10456, LDPC_TABLE_DATA_WIDTH)),
    4016 => std_logic_vector(to_unsigned(9774, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4017 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4018 => std_logic_vector(to_unsigned(1692, LDPC_TABLE_DATA_WIDTH)),
    4019 => std_logic_vector(to_unsigned(9276, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4020 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4021 => std_logic_vector(to_unsigned(10037, LDPC_TABLE_DATA_WIDTH)),
    4022 => std_logic_vector(to_unsigned(4038, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4023 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4024 => std_logic_vector(to_unsigned(3964, LDPC_TABLE_DATA_WIDTH)),
    4025 => std_logic_vector(to_unsigned(338, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4026 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4027 => std_logic_vector(to_unsigned(2640, LDPC_TABLE_DATA_WIDTH)),
    4028 => std_logic_vector(to_unsigned(5087, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4029 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4030 => std_logic_vector(to_unsigned(858, LDPC_TABLE_DATA_WIDTH)),
    4031 => std_logic_vector(to_unsigned(3473, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4032 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4033 => std_logic_vector(to_unsigned(5582, LDPC_TABLE_DATA_WIDTH)),
    4034 => std_logic_vector(to_unsigned(5683, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4035 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4036 => std_logic_vector(to_unsigned(9523, LDPC_TABLE_DATA_WIDTH)),
    4037 => std_logic_vector(to_unsigned(916, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4038 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4039 => std_logic_vector(to_unsigned(4107, LDPC_TABLE_DATA_WIDTH)),
    4040 => std_logic_vector(to_unsigned(1559, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4041 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4042 => std_logic_vector(to_unsigned(4506, LDPC_TABLE_DATA_WIDTH)),
    4043 => std_logic_vector(to_unsigned(3491, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4044 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4045 => std_logic_vector(to_unsigned(8191, LDPC_TABLE_DATA_WIDTH)),
    4046 => std_logic_vector(to_unsigned(4182, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4047 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4048 => std_logic_vector(to_unsigned(10192, LDPC_TABLE_DATA_WIDTH)),
    4049 => std_logic_vector(to_unsigned(6157, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4050 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4051 => std_logic_vector(to_unsigned(5668, LDPC_TABLE_DATA_WIDTH)),
    4052 => std_logic_vector(to_unsigned(3305, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4053 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4054 => std_logic_vector(to_unsigned(3449, LDPC_TABLE_DATA_WIDTH)),
    4055 => std_logic_vector(to_unsigned(1540, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4056 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    4057 => std_logic_vector(to_unsigned(4766, LDPC_TABLE_DATA_WIDTH)),
    4058 => std_logic_vector(to_unsigned(2697, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4059 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    4060 => std_logic_vector(to_unsigned(4069, LDPC_TABLE_DATA_WIDTH)),
    4061 => std_logic_vector(to_unsigned(6675, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4062 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    4063 => std_logic_vector(to_unsigned(1117, LDPC_TABLE_DATA_WIDTH)),
    4064 => std_logic_vector(to_unsigned(1016, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4065 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    4066 => std_logic_vector(to_unsigned(5619, LDPC_TABLE_DATA_WIDTH)),
    4067 => std_logic_vector(to_unsigned(3085, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4068 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    4069 => std_logic_vector(to_unsigned(8483, LDPC_TABLE_DATA_WIDTH)),
    4070 => std_logic_vector(to_unsigned(8400, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4071 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    4072 => std_logic_vector(to_unsigned(8255, LDPC_TABLE_DATA_WIDTH)),
    4073 => std_logic_vector(to_unsigned(394, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4074 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    4075 => std_logic_vector(to_unsigned(6338, LDPC_TABLE_DATA_WIDTH)),
    4076 => std_logic_vector(to_unsigned(5042, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4077 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    4078 => std_logic_vector(to_unsigned(6174, LDPC_TABLE_DATA_WIDTH)),
    4079 => std_logic_vector(to_unsigned(5119, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4080 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    4081 => std_logic_vector(to_unsigned(7203, LDPC_TABLE_DATA_WIDTH)),
    4082 => std_logic_vector(to_unsigned(1989, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4083 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    4084 => std_logic_vector(to_unsigned(1781, LDPC_TABLE_DATA_WIDTH)),
    4085 => std_logic_vector(to_unsigned(5174, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4086 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4087 => std_logic_vector(to_unsigned(1464, LDPC_TABLE_DATA_WIDTH)),
    4088 => std_logic_vector(to_unsigned(3559, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4089 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4090 => std_logic_vector(to_unsigned(3376, LDPC_TABLE_DATA_WIDTH)),
    4091 => std_logic_vector(to_unsigned(4214, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4092 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4093 => std_logic_vector(to_unsigned(7238, LDPC_TABLE_DATA_WIDTH)),
    4094 => std_logic_vector(to_unsigned(67, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4095 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4096 => std_logic_vector(to_unsigned(10595, LDPC_TABLE_DATA_WIDTH)),
    4097 => std_logic_vector(to_unsigned(8831, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4098 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4099 => std_logic_vector(to_unsigned(1221, LDPC_TABLE_DATA_WIDTH)),
    4100 => std_logic_vector(to_unsigned(6513, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4101 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4102 => std_logic_vector(to_unsigned(5300, LDPC_TABLE_DATA_WIDTH)),
    4103 => std_logic_vector(to_unsigned(4652, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4104 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4105 => std_logic_vector(to_unsigned(1429, LDPC_TABLE_DATA_WIDTH)),
    4106 => std_logic_vector(to_unsigned(9749, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4107 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4108 => std_logic_vector(to_unsigned(7878, LDPC_TABLE_DATA_WIDTH)),
    4109 => std_logic_vector(to_unsigned(5131, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4110 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4111 => std_logic_vector(to_unsigned(4435, LDPC_TABLE_DATA_WIDTH)),
    4112 => std_logic_vector(to_unsigned(10284, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4113 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4114 => std_logic_vector(to_unsigned(6331, LDPC_TABLE_DATA_WIDTH)),
    4115 => std_logic_vector(to_unsigned(5507, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4116 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4117 => std_logic_vector(to_unsigned(6662, LDPC_TABLE_DATA_WIDTH)),
    4118 => std_logic_vector(to_unsigned(4941, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4119 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4120 => std_logic_vector(to_unsigned(9614, LDPC_TABLE_DATA_WIDTH)),
    4121 => std_logic_vector(to_unsigned(10238, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4122 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4123 => std_logic_vector(to_unsigned(8400, LDPC_TABLE_DATA_WIDTH)),
    4124 => std_logic_vector(to_unsigned(8025, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4125 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4126 => std_logic_vector(to_unsigned(9156, LDPC_TABLE_DATA_WIDTH)),
    4127 => std_logic_vector(to_unsigned(5630, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4128 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4129 => std_logic_vector(to_unsigned(7067, LDPC_TABLE_DATA_WIDTH)),
    4130 => std_logic_vector(to_unsigned(8878, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4131 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4132 => std_logic_vector(to_unsigned(9027, LDPC_TABLE_DATA_WIDTH)),
    4133 => std_logic_vector(to_unsigned(3415, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4134 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4135 => std_logic_vector(to_unsigned(1690, LDPC_TABLE_DATA_WIDTH)),
    4136 => std_logic_vector(to_unsigned(3866, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4137 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4138 => std_logic_vector(to_unsigned(2854, LDPC_TABLE_DATA_WIDTH)),
    4139 => std_logic_vector(to_unsigned(8469, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4140 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4141 => std_logic_vector(to_unsigned(6206, LDPC_TABLE_DATA_WIDTH)),
    4142 => std_logic_vector(to_unsigned(630, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4143 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4144 => std_logic_vector(to_unsigned(363, LDPC_TABLE_DATA_WIDTH)),
    4145 => std_logic_vector(to_unsigned(5453, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4146 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    4147 => std_logic_vector(to_unsigned(4125, LDPC_TABLE_DATA_WIDTH)),
    4148 => std_logic_vector(to_unsigned(7008, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4149 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    4150 => std_logic_vector(to_unsigned(1612, LDPC_TABLE_DATA_WIDTH)),
    4151 => std_logic_vector(to_unsigned(6702, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4152 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    4153 => std_logic_vector(to_unsigned(9069, LDPC_TABLE_DATA_WIDTH)),
    4154 => std_logic_vector(to_unsigned(9226, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4155 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    4156 => std_logic_vector(to_unsigned(5767, LDPC_TABLE_DATA_WIDTH)),
    4157 => std_logic_vector(to_unsigned(4060, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4158 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    4159 => std_logic_vector(to_unsigned(3743, LDPC_TABLE_DATA_WIDTH)),
    4160 => std_logic_vector(to_unsigned(9237, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4161 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    4162 => std_logic_vector(to_unsigned(7018, LDPC_TABLE_DATA_WIDTH)),
    4163 => std_logic_vector(to_unsigned(5572, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4164 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    4165 => std_logic_vector(to_unsigned(8892, LDPC_TABLE_DATA_WIDTH)),
    4166 => std_logic_vector(to_unsigned(4536, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4167 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    4168 => std_logic_vector(to_unsigned(853, LDPC_TABLE_DATA_WIDTH)),
    4169 => std_logic_vector(to_unsigned(6064, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4170 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    4171 => std_logic_vector(to_unsigned(8069, LDPC_TABLE_DATA_WIDTH)),
    4172 => std_logic_vector(to_unsigned(5893, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4173 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    4174 => std_logic_vector(to_unsigned(2051, LDPC_TABLE_DATA_WIDTH)),
    4175 => std_logic_vector(to_unsigned(2885, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4176 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4177 => std_logic_vector(to_unsigned(10691, LDPC_TABLE_DATA_WIDTH)),
    4178 => std_logic_vector(to_unsigned(3153, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4179 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4180 => std_logic_vector(to_unsigned(3602, LDPC_TABLE_DATA_WIDTH)),
    4181 => std_logic_vector(to_unsigned(4055, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4182 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4183 => std_logic_vector(to_unsigned(328, LDPC_TABLE_DATA_WIDTH)),
    4184 => std_logic_vector(to_unsigned(1717, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4185 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4186 => std_logic_vector(to_unsigned(2219, LDPC_TABLE_DATA_WIDTH)),
    4187 => std_logic_vector(to_unsigned(9299, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4188 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4189 => std_logic_vector(to_unsigned(1939, LDPC_TABLE_DATA_WIDTH)),
    4190 => std_logic_vector(to_unsigned(7898, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4191 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4192 => std_logic_vector(to_unsigned(617, LDPC_TABLE_DATA_WIDTH)),
    4193 => std_logic_vector(to_unsigned(206, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4194 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4195 => std_logic_vector(to_unsigned(8544, LDPC_TABLE_DATA_WIDTH)),
    4196 => std_logic_vector(to_unsigned(1374, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4197 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4198 => std_logic_vector(to_unsigned(10676, LDPC_TABLE_DATA_WIDTH)),
    4199 => std_logic_vector(to_unsigned(3240, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4200 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4201 => std_logic_vector(to_unsigned(6672, LDPC_TABLE_DATA_WIDTH)),
    4202 => std_logic_vector(to_unsigned(9489, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4203 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4204 => std_logic_vector(to_unsigned(3170, LDPC_TABLE_DATA_WIDTH)),
    4205 => std_logic_vector(to_unsigned(7457, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4206 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4207 => std_logic_vector(to_unsigned(7868, LDPC_TABLE_DATA_WIDTH)),
    4208 => std_logic_vector(to_unsigned(5731, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4209 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4210 => std_logic_vector(to_unsigned(6121, LDPC_TABLE_DATA_WIDTH)),
    4211 => std_logic_vector(to_unsigned(10732, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4212 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4213 => std_logic_vector(to_unsigned(4843, LDPC_TABLE_DATA_WIDTH)),
    4214 => std_logic_vector(to_unsigned(9132, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4215 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4216 => std_logic_vector(to_unsigned(580, LDPC_TABLE_DATA_WIDTH)),
    4217 => std_logic_vector(to_unsigned(9591, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4218 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4219 => std_logic_vector(to_unsigned(6267, LDPC_TABLE_DATA_WIDTH)),
    4220 => std_logic_vector(to_unsigned(9290, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4221 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4222 => std_logic_vector(to_unsigned(3009, LDPC_TABLE_DATA_WIDTH)),
    4223 => std_logic_vector(to_unsigned(2268, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4224 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4225 => std_logic_vector(to_unsigned(195, LDPC_TABLE_DATA_WIDTH)),
    4226 => std_logic_vector(to_unsigned(2419, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4227 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4228 => std_logic_vector(to_unsigned(8016, LDPC_TABLE_DATA_WIDTH)),
    4229 => std_logic_vector(to_unsigned(1557, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4230 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4231 => std_logic_vector(to_unsigned(1516, LDPC_TABLE_DATA_WIDTH)),
    4232 => std_logic_vector(to_unsigned(9195, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4233 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4234 => std_logic_vector(to_unsigned(8062, LDPC_TABLE_DATA_WIDTH)),
    4235 => std_logic_vector(to_unsigned(9064, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4236 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    4237 => std_logic_vector(to_unsigned(2095, LDPC_TABLE_DATA_WIDTH)),
    4238 => std_logic_vector(to_unsigned(8968, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4239 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    4240 => std_logic_vector(to_unsigned(753, LDPC_TABLE_DATA_WIDTH)),
    4241 => std_logic_vector(to_unsigned(7326, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4242 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    4243 => std_logic_vector(to_unsigned(6291, LDPC_TABLE_DATA_WIDTH)),
    4244 => std_logic_vector(to_unsigned(3833, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4245 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    4246 => std_logic_vector(to_unsigned(2614, LDPC_TABLE_DATA_WIDTH)),
    4247 => std_logic_vector(to_unsigned(7844, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4248 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    4249 => std_logic_vector(to_unsigned(2303, LDPC_TABLE_DATA_WIDTH)),
    4250 => std_logic_vector(to_unsigned(646, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4251 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    4252 => std_logic_vector(to_unsigned(2075, LDPC_TABLE_DATA_WIDTH)),
    4253 => std_logic_vector(to_unsigned(611, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4254 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    4255 => std_logic_vector(to_unsigned(4687, LDPC_TABLE_DATA_WIDTH)),
    4256 => std_logic_vector(to_unsigned(362, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4257 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    4258 => std_logic_vector(to_unsigned(8684, LDPC_TABLE_DATA_WIDTH)),
    4259 => std_logic_vector(to_unsigned(9940, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4260 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    4261 => std_logic_vector(to_unsigned(4830, LDPC_TABLE_DATA_WIDTH)),
    4262 => std_logic_vector(to_unsigned(2065, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4263 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    4264 => std_logic_vector(to_unsigned(7038, LDPC_TABLE_DATA_WIDTH)),
    4265 => std_logic_vector(to_unsigned(1363, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4266 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4267 => std_logic_vector(to_unsigned(1769, LDPC_TABLE_DATA_WIDTH)),
    4268 => std_logic_vector(to_unsigned(7837, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4269 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4270 => std_logic_vector(to_unsigned(3801, LDPC_TABLE_DATA_WIDTH)),
    4271 => std_logic_vector(to_unsigned(1689, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4272 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4273 => std_logic_vector(to_unsigned(10070, LDPC_TABLE_DATA_WIDTH)),
    4274 => std_logic_vector(to_unsigned(2359, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4275 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4276 => std_logic_vector(to_unsigned(3667, LDPC_TABLE_DATA_WIDTH)),
    4277 => std_logic_vector(to_unsigned(9918, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4278 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4279 => std_logic_vector(to_unsigned(1914, LDPC_TABLE_DATA_WIDTH)),
    4280 => std_logic_vector(to_unsigned(6920, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4281 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4282 => std_logic_vector(to_unsigned(4244, LDPC_TABLE_DATA_WIDTH)),
    4283 => std_logic_vector(to_unsigned(5669, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4284 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4285 => std_logic_vector(to_unsigned(10245, LDPC_TABLE_DATA_WIDTH)),
    4286 => std_logic_vector(to_unsigned(7821, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4287 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4288 => std_logic_vector(to_unsigned(7648, LDPC_TABLE_DATA_WIDTH)),
    4289 => std_logic_vector(to_unsigned(3944, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4290 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4291 => std_logic_vector(to_unsigned(3310, LDPC_TABLE_DATA_WIDTH)),
    4292 => std_logic_vector(to_unsigned(5488, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4293 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4294 => std_logic_vector(to_unsigned(6346, LDPC_TABLE_DATA_WIDTH)),
    4295 => std_logic_vector(to_unsigned(9666, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4296 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4297 => std_logic_vector(to_unsigned(7088, LDPC_TABLE_DATA_WIDTH)),
    4298 => std_logic_vector(to_unsigned(6122, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4299 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4300 => std_logic_vector(to_unsigned(1291, LDPC_TABLE_DATA_WIDTH)),
    4301 => std_logic_vector(to_unsigned(7827, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4302 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4303 => std_logic_vector(to_unsigned(10592, LDPC_TABLE_DATA_WIDTH)),
    4304 => std_logic_vector(to_unsigned(8945, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4305 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4306 => std_logic_vector(to_unsigned(3609, LDPC_TABLE_DATA_WIDTH)),
    4307 => std_logic_vector(to_unsigned(7120, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4308 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4309 => std_logic_vector(to_unsigned(9168, LDPC_TABLE_DATA_WIDTH)),
    4310 => std_logic_vector(to_unsigned(9112, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4311 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4312 => std_logic_vector(to_unsigned(6203, LDPC_TABLE_DATA_WIDTH)),
    4313 => std_logic_vector(to_unsigned(8052, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4314 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4315 => std_logic_vector(to_unsigned(3330, LDPC_TABLE_DATA_WIDTH)),
    4316 => std_logic_vector(to_unsigned(2895, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4317 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4318 => std_logic_vector(to_unsigned(4264, LDPC_TABLE_DATA_WIDTH)),
    4319 => std_logic_vector(to_unsigned(10563, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4320 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4321 => std_logic_vector(to_unsigned(10556, LDPC_TABLE_DATA_WIDTH)),
    4322 => std_logic_vector(to_unsigned(6496, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4323 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4324 => std_logic_vector(to_unsigned(8807, LDPC_TABLE_DATA_WIDTH)),
    4325 => std_logic_vector(to_unsigned(7645, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4326 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    4327 => std_logic_vector(to_unsigned(1999, LDPC_TABLE_DATA_WIDTH)),
    4328 => std_logic_vector(to_unsigned(4530, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4329 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    4330 => std_logic_vector(to_unsigned(9202, LDPC_TABLE_DATA_WIDTH)),
    4331 => std_logic_vector(to_unsigned(6818, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4332 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    4333 => std_logic_vector(to_unsigned(3403, LDPC_TABLE_DATA_WIDTH)),
    4334 => std_logic_vector(to_unsigned(1734, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4335 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    4336 => std_logic_vector(to_unsigned(2106, LDPC_TABLE_DATA_WIDTH)),
    4337 => std_logic_vector(to_unsigned(9023, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4338 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    4339 => std_logic_vector(to_unsigned(6881, LDPC_TABLE_DATA_WIDTH)),
    4340 => std_logic_vector(to_unsigned(3883, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4341 => std_logic_vector(to_unsigned(25, LDPC_TABLE_DATA_WIDTH)),
    4342 => std_logic_vector(to_unsigned(3895, LDPC_TABLE_DATA_WIDTH)),
    4343 => std_logic_vector(to_unsigned(2171, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4344 => std_logic_vector(to_unsigned(26, LDPC_TABLE_DATA_WIDTH)),
    4345 => std_logic_vector(to_unsigned(4062, LDPC_TABLE_DATA_WIDTH)),
    4346 => std_logic_vector(to_unsigned(6424, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4347 => std_logic_vector(to_unsigned(27, LDPC_TABLE_DATA_WIDTH)),
    4348 => std_logic_vector(to_unsigned(3755, LDPC_TABLE_DATA_WIDTH)),
    4349 => std_logic_vector(to_unsigned(9536, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4350 => std_logic_vector(to_unsigned(28, LDPC_TABLE_DATA_WIDTH)),
    4351 => std_logic_vector(to_unsigned(4683, LDPC_TABLE_DATA_WIDTH)),
    4352 => std_logic_vector(to_unsigned(2131, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4353 => std_logic_vector(to_unsigned(29, LDPC_TABLE_DATA_WIDTH)),
    4354 => std_logic_vector(to_unsigned(7347, LDPC_TABLE_DATA_WIDTH)),
    4355 => std_logic_vector(to_unsigned(8027, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C8_9
    4356 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4357 => std_logic_vector(to_unsigned(6235, LDPC_TABLE_DATA_WIDTH)),
    4358 => std_logic_vector(to_unsigned(2848, LDPC_TABLE_DATA_WIDTH)),
    4359 => std_logic_vector(to_unsigned(3222, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4360 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4361 => std_logic_vector(to_unsigned(5800, LDPC_TABLE_DATA_WIDTH)),
    4362 => std_logic_vector(to_unsigned(3492, LDPC_TABLE_DATA_WIDTH)),
    4363 => std_logic_vector(to_unsigned(5348, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4364 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4365 => std_logic_vector(to_unsigned(2757, LDPC_TABLE_DATA_WIDTH)),
    4366 => std_logic_vector(to_unsigned(927, LDPC_TABLE_DATA_WIDTH)),
    4367 => std_logic_vector(to_unsigned(90, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4368 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4369 => std_logic_vector(to_unsigned(6961, LDPC_TABLE_DATA_WIDTH)),
    4370 => std_logic_vector(to_unsigned(4516, LDPC_TABLE_DATA_WIDTH)),
    4371 => std_logic_vector(to_unsigned(4739, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4372 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4373 => std_logic_vector(to_unsigned(1172, LDPC_TABLE_DATA_WIDTH)),
    4374 => std_logic_vector(to_unsigned(3237, LDPC_TABLE_DATA_WIDTH)),
    4375 => std_logic_vector(to_unsigned(6264, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4376 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4377 => std_logic_vector(to_unsigned(1927, LDPC_TABLE_DATA_WIDTH)),
    4378 => std_logic_vector(to_unsigned(2425, LDPC_TABLE_DATA_WIDTH)),
    4379 => std_logic_vector(to_unsigned(3683, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4380 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4381 => std_logic_vector(to_unsigned(3714, LDPC_TABLE_DATA_WIDTH)),
    4382 => std_logic_vector(to_unsigned(6309, LDPC_TABLE_DATA_WIDTH)),
    4383 => std_logic_vector(to_unsigned(2495, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4384 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4385 => std_logic_vector(to_unsigned(3070, LDPC_TABLE_DATA_WIDTH)),
    4386 => std_logic_vector(to_unsigned(6342, LDPC_TABLE_DATA_WIDTH)),
    4387 => std_logic_vector(to_unsigned(7154, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4388 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4389 => std_logic_vector(to_unsigned(2428, LDPC_TABLE_DATA_WIDTH)),
    4390 => std_logic_vector(to_unsigned(613, LDPC_TABLE_DATA_WIDTH)),
    4391 => std_logic_vector(to_unsigned(3761, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4392 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4393 => std_logic_vector(to_unsigned(2906, LDPC_TABLE_DATA_WIDTH)),
    4394 => std_logic_vector(to_unsigned(264, LDPC_TABLE_DATA_WIDTH)),
    4395 => std_logic_vector(to_unsigned(5927, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4396 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4397 => std_logic_vector(to_unsigned(1716, LDPC_TABLE_DATA_WIDTH)),
    4398 => std_logic_vector(to_unsigned(1950, LDPC_TABLE_DATA_WIDTH)),
    4399 => std_logic_vector(to_unsigned(4273, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4400 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4401 => std_logic_vector(to_unsigned(4613, LDPC_TABLE_DATA_WIDTH)),
    4402 => std_logic_vector(to_unsigned(6179, LDPC_TABLE_DATA_WIDTH)),
    4403 => std_logic_vector(to_unsigned(3491, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4404 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4405 => std_logic_vector(to_unsigned(4865, LDPC_TABLE_DATA_WIDTH)),
    4406 => std_logic_vector(to_unsigned(3286, LDPC_TABLE_DATA_WIDTH)),
    4407 => std_logic_vector(to_unsigned(6005, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4408 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4409 => std_logic_vector(to_unsigned(1343, LDPC_TABLE_DATA_WIDTH)),
    4410 => std_logic_vector(to_unsigned(5923, LDPC_TABLE_DATA_WIDTH)),
    4411 => std_logic_vector(to_unsigned(3529, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4412 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4413 => std_logic_vector(to_unsigned(4589, LDPC_TABLE_DATA_WIDTH)),
    4414 => std_logic_vector(to_unsigned(4035, LDPC_TABLE_DATA_WIDTH)),
    4415 => std_logic_vector(to_unsigned(2132, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4416 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4417 => std_logic_vector(to_unsigned(1579, LDPC_TABLE_DATA_WIDTH)),
    4418 => std_logic_vector(to_unsigned(3920, LDPC_TABLE_DATA_WIDTH)),
    4419 => std_logic_vector(to_unsigned(6737, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4420 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4421 => std_logic_vector(to_unsigned(1644, LDPC_TABLE_DATA_WIDTH)),
    4422 => std_logic_vector(to_unsigned(1191, LDPC_TABLE_DATA_WIDTH)),
    4423 => std_logic_vector(to_unsigned(5998, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4424 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4425 => std_logic_vector(to_unsigned(1482, LDPC_TABLE_DATA_WIDTH)),
    4426 => std_logic_vector(to_unsigned(2381, LDPC_TABLE_DATA_WIDTH)),
    4427 => std_logic_vector(to_unsigned(4620, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4428 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4429 => std_logic_vector(to_unsigned(6791, LDPC_TABLE_DATA_WIDTH)),
    4430 => std_logic_vector(to_unsigned(6014, LDPC_TABLE_DATA_WIDTH)),
    4431 => std_logic_vector(to_unsigned(6596, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4432 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4433 => std_logic_vector(to_unsigned(2738, LDPC_TABLE_DATA_WIDTH)),
    4434 => std_logic_vector(to_unsigned(5918, LDPC_TABLE_DATA_WIDTH)),
    4435 => std_logic_vector(to_unsigned(3786, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4436 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4437 => std_logic_vector(to_unsigned(5156, LDPC_TABLE_DATA_WIDTH)),
    4438 => std_logic_vector(to_unsigned(6166, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4439 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4440 => std_logic_vector(to_unsigned(1504, LDPC_TABLE_DATA_WIDTH)),
    4441 => std_logic_vector(to_unsigned(4356, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4442 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4443 => std_logic_vector(to_unsigned(130, LDPC_TABLE_DATA_WIDTH)),
    4444 => std_logic_vector(to_unsigned(1904, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4445 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4446 => std_logic_vector(to_unsigned(6027, LDPC_TABLE_DATA_WIDTH)),
    4447 => std_logic_vector(to_unsigned(3187, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4448 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4449 => std_logic_vector(to_unsigned(6718, LDPC_TABLE_DATA_WIDTH)),
    4450 => std_logic_vector(to_unsigned(759, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4451 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4452 => std_logic_vector(to_unsigned(6240, LDPC_TABLE_DATA_WIDTH)),
    4453 => std_logic_vector(to_unsigned(2870, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4454 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4455 => std_logic_vector(to_unsigned(2343, LDPC_TABLE_DATA_WIDTH)),
    4456 => std_logic_vector(to_unsigned(1311, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4457 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4458 => std_logic_vector(to_unsigned(1039, LDPC_TABLE_DATA_WIDTH)),
    4459 => std_logic_vector(to_unsigned(5465, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4460 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4461 => std_logic_vector(to_unsigned(6617, LDPC_TABLE_DATA_WIDTH)),
    4462 => std_logic_vector(to_unsigned(2513, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4463 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4464 => std_logic_vector(to_unsigned(1588, LDPC_TABLE_DATA_WIDTH)),
    4465 => std_logic_vector(to_unsigned(5222, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4466 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4467 => std_logic_vector(to_unsigned(6561, LDPC_TABLE_DATA_WIDTH)),
    4468 => std_logic_vector(to_unsigned(535, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4469 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4470 => std_logic_vector(to_unsigned(4765, LDPC_TABLE_DATA_WIDTH)),
    4471 => std_logic_vector(to_unsigned(2054, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4472 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4473 => std_logic_vector(to_unsigned(5966, LDPC_TABLE_DATA_WIDTH)),
    4474 => std_logic_vector(to_unsigned(6892, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4475 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4476 => std_logic_vector(to_unsigned(1969, LDPC_TABLE_DATA_WIDTH)),
    4477 => std_logic_vector(to_unsigned(3869, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4478 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4479 => std_logic_vector(to_unsigned(3571, LDPC_TABLE_DATA_WIDTH)),
    4480 => std_logic_vector(to_unsigned(2420, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4481 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4482 => std_logic_vector(to_unsigned(4632, LDPC_TABLE_DATA_WIDTH)),
    4483 => std_logic_vector(to_unsigned(981, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4484 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4485 => std_logic_vector(to_unsigned(3215, LDPC_TABLE_DATA_WIDTH)),
    4486 => std_logic_vector(to_unsigned(4163, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4487 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4488 => std_logic_vector(to_unsigned(973, LDPC_TABLE_DATA_WIDTH)),
    4489 => std_logic_vector(to_unsigned(3117, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4490 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4491 => std_logic_vector(to_unsigned(3802, LDPC_TABLE_DATA_WIDTH)),
    4492 => std_logic_vector(to_unsigned(6198, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4493 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4494 => std_logic_vector(to_unsigned(3794, LDPC_TABLE_DATA_WIDTH)),
    4495 => std_logic_vector(to_unsigned(3948, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4496 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4497 => std_logic_vector(to_unsigned(3196, LDPC_TABLE_DATA_WIDTH)),
    4498 => std_logic_vector(to_unsigned(6126, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4499 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4500 => std_logic_vector(to_unsigned(573, LDPC_TABLE_DATA_WIDTH)),
    4501 => std_logic_vector(to_unsigned(1909, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4502 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4503 => std_logic_vector(to_unsigned(850, LDPC_TABLE_DATA_WIDTH)),
    4504 => std_logic_vector(to_unsigned(4034, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4505 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4506 => std_logic_vector(to_unsigned(5622, LDPC_TABLE_DATA_WIDTH)),
    4507 => std_logic_vector(to_unsigned(1601, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4508 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4509 => std_logic_vector(to_unsigned(6005, LDPC_TABLE_DATA_WIDTH)),
    4510 => std_logic_vector(to_unsigned(524, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4511 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4512 => std_logic_vector(to_unsigned(5251, LDPC_TABLE_DATA_WIDTH)),
    4513 => std_logic_vector(to_unsigned(5783, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4514 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4515 => std_logic_vector(to_unsigned(172, LDPC_TABLE_DATA_WIDTH)),
    4516 => std_logic_vector(to_unsigned(2032, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4517 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4518 => std_logic_vector(to_unsigned(1875, LDPC_TABLE_DATA_WIDTH)),
    4519 => std_logic_vector(to_unsigned(2475, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4520 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4521 => std_logic_vector(to_unsigned(497, LDPC_TABLE_DATA_WIDTH)),
    4522 => std_logic_vector(to_unsigned(1291, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4523 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4524 => std_logic_vector(to_unsigned(2566, LDPC_TABLE_DATA_WIDTH)),
    4525 => std_logic_vector(to_unsigned(3430, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4526 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4527 => std_logic_vector(to_unsigned(1249, LDPC_TABLE_DATA_WIDTH)),
    4528 => std_logic_vector(to_unsigned(740, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4529 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4530 => std_logic_vector(to_unsigned(2944, LDPC_TABLE_DATA_WIDTH)),
    4531 => std_logic_vector(to_unsigned(1948, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4532 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4533 => std_logic_vector(to_unsigned(6528, LDPC_TABLE_DATA_WIDTH)),
    4534 => std_logic_vector(to_unsigned(2899, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4535 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4536 => std_logic_vector(to_unsigned(2243, LDPC_TABLE_DATA_WIDTH)),
    4537 => std_logic_vector(to_unsigned(3616, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4538 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4539 => std_logic_vector(to_unsigned(867, LDPC_TABLE_DATA_WIDTH)),
    4540 => std_logic_vector(to_unsigned(3733, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4541 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4542 => std_logic_vector(to_unsigned(1374, LDPC_TABLE_DATA_WIDTH)),
    4543 => std_logic_vector(to_unsigned(4702, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4544 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4545 => std_logic_vector(to_unsigned(4698, LDPC_TABLE_DATA_WIDTH)),
    4546 => std_logic_vector(to_unsigned(2285, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4547 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4548 => std_logic_vector(to_unsigned(4760, LDPC_TABLE_DATA_WIDTH)),
    4549 => std_logic_vector(to_unsigned(3917, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4550 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4551 => std_logic_vector(to_unsigned(1859, LDPC_TABLE_DATA_WIDTH)),
    4552 => std_logic_vector(to_unsigned(4058, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4553 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4554 => std_logic_vector(to_unsigned(6141, LDPC_TABLE_DATA_WIDTH)),
    4555 => std_logic_vector(to_unsigned(3527, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4556 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4557 => std_logic_vector(to_unsigned(2148, LDPC_TABLE_DATA_WIDTH)),
    4558 => std_logic_vector(to_unsigned(5066, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4559 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4560 => std_logic_vector(to_unsigned(1306, LDPC_TABLE_DATA_WIDTH)),
    4561 => std_logic_vector(to_unsigned(145, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4562 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4563 => std_logic_vector(to_unsigned(2319, LDPC_TABLE_DATA_WIDTH)),
    4564 => std_logic_vector(to_unsigned(871, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4565 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4566 => std_logic_vector(to_unsigned(3463, LDPC_TABLE_DATA_WIDTH)),
    4567 => std_logic_vector(to_unsigned(1061, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4568 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4569 => std_logic_vector(to_unsigned(5554, LDPC_TABLE_DATA_WIDTH)),
    4570 => std_logic_vector(to_unsigned(6647, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4571 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4572 => std_logic_vector(to_unsigned(5837, LDPC_TABLE_DATA_WIDTH)),
    4573 => std_logic_vector(to_unsigned(339, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4574 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4575 => std_logic_vector(to_unsigned(5821, LDPC_TABLE_DATA_WIDTH)),
    4576 => std_logic_vector(to_unsigned(4932, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4577 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4578 => std_logic_vector(to_unsigned(6356, LDPC_TABLE_DATA_WIDTH)),
    4579 => std_logic_vector(to_unsigned(4756, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4580 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4581 => std_logic_vector(to_unsigned(3930, LDPC_TABLE_DATA_WIDTH)),
    4582 => std_logic_vector(to_unsigned(418, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4583 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4584 => std_logic_vector(to_unsigned(211, LDPC_TABLE_DATA_WIDTH)),
    4585 => std_logic_vector(to_unsigned(3094, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4586 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4587 => std_logic_vector(to_unsigned(1007, LDPC_TABLE_DATA_WIDTH)),
    4588 => std_logic_vector(to_unsigned(4928, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4589 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4590 => std_logic_vector(to_unsigned(3584, LDPC_TABLE_DATA_WIDTH)),
    4591 => std_logic_vector(to_unsigned(1235, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4592 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4593 => std_logic_vector(to_unsigned(6982, LDPC_TABLE_DATA_WIDTH)),
    4594 => std_logic_vector(to_unsigned(2869, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4595 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4596 => std_logic_vector(to_unsigned(1612, LDPC_TABLE_DATA_WIDTH)),
    4597 => std_logic_vector(to_unsigned(1013, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4598 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4599 => std_logic_vector(to_unsigned(953, LDPC_TABLE_DATA_WIDTH)),
    4600 => std_logic_vector(to_unsigned(4964, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4601 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4602 => std_logic_vector(to_unsigned(4555, LDPC_TABLE_DATA_WIDTH)),
    4603 => std_logic_vector(to_unsigned(4410, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4604 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4605 => std_logic_vector(to_unsigned(4925, LDPC_TABLE_DATA_WIDTH)),
    4606 => std_logic_vector(to_unsigned(4842, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4607 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4608 => std_logic_vector(to_unsigned(5778, LDPC_TABLE_DATA_WIDTH)),
    4609 => std_logic_vector(to_unsigned(600, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4610 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4611 => std_logic_vector(to_unsigned(6509, LDPC_TABLE_DATA_WIDTH)),
    4612 => std_logic_vector(to_unsigned(2417, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4613 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4614 => std_logic_vector(to_unsigned(1260, LDPC_TABLE_DATA_WIDTH)),
    4615 => std_logic_vector(to_unsigned(4903, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4616 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4617 => std_logic_vector(to_unsigned(3369, LDPC_TABLE_DATA_WIDTH)),
    4618 => std_logic_vector(to_unsigned(3031, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4619 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4620 => std_logic_vector(to_unsigned(3557, LDPC_TABLE_DATA_WIDTH)),
    4621 => std_logic_vector(to_unsigned(3224, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4622 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4623 => std_logic_vector(to_unsigned(3028, LDPC_TABLE_DATA_WIDTH)),
    4624 => std_logic_vector(to_unsigned(583, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4625 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4626 => std_logic_vector(to_unsigned(3258, LDPC_TABLE_DATA_WIDTH)),
    4627 => std_logic_vector(to_unsigned(440, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4628 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4629 => std_logic_vector(to_unsigned(6226, LDPC_TABLE_DATA_WIDTH)),
    4630 => std_logic_vector(to_unsigned(6655, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4631 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4632 => std_logic_vector(to_unsigned(4895, LDPC_TABLE_DATA_WIDTH)),
    4633 => std_logic_vector(to_unsigned(1094, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4634 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4635 => std_logic_vector(to_unsigned(1481, LDPC_TABLE_DATA_WIDTH)),
    4636 => std_logic_vector(to_unsigned(6847, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4637 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4638 => std_logic_vector(to_unsigned(4433, LDPC_TABLE_DATA_WIDTH)),
    4639 => std_logic_vector(to_unsigned(1932, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4640 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4641 => std_logic_vector(to_unsigned(2107, LDPC_TABLE_DATA_WIDTH)),
    4642 => std_logic_vector(to_unsigned(1649, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4643 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4644 => std_logic_vector(to_unsigned(2119, LDPC_TABLE_DATA_WIDTH)),
    4645 => std_logic_vector(to_unsigned(2065, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4646 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4647 => std_logic_vector(to_unsigned(4003, LDPC_TABLE_DATA_WIDTH)),
    4648 => std_logic_vector(to_unsigned(6388, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4649 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4650 => std_logic_vector(to_unsigned(6720, LDPC_TABLE_DATA_WIDTH)),
    4651 => std_logic_vector(to_unsigned(3622, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4652 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4653 => std_logic_vector(to_unsigned(3694, LDPC_TABLE_DATA_WIDTH)),
    4654 => std_logic_vector(to_unsigned(4521, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4655 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4656 => std_logic_vector(to_unsigned(1164, LDPC_TABLE_DATA_WIDTH)),
    4657 => std_logic_vector(to_unsigned(7050, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4658 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4659 => std_logic_vector(to_unsigned(1965, LDPC_TABLE_DATA_WIDTH)),
    4660 => std_logic_vector(to_unsigned(3613, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4661 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4662 => std_logic_vector(to_unsigned(4331, LDPC_TABLE_DATA_WIDTH)),
    4663 => std_logic_vector(to_unsigned(66, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4664 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4665 => std_logic_vector(to_unsigned(2970, LDPC_TABLE_DATA_WIDTH)),
    4666 => std_logic_vector(to_unsigned(1796, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4667 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4668 => std_logic_vector(to_unsigned(4652, LDPC_TABLE_DATA_WIDTH)),
    4669 => std_logic_vector(to_unsigned(3218, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4670 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4671 => std_logic_vector(to_unsigned(1762, LDPC_TABLE_DATA_WIDTH)),
    4672 => std_logic_vector(to_unsigned(4777, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4673 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4674 => std_logic_vector(to_unsigned(5736, LDPC_TABLE_DATA_WIDTH)),
    4675 => std_logic_vector(to_unsigned(1399, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4676 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4677 => std_logic_vector(to_unsigned(970, LDPC_TABLE_DATA_WIDTH)),
    4678 => std_logic_vector(to_unsigned(2572, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4679 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4680 => std_logic_vector(to_unsigned(2062, LDPC_TABLE_DATA_WIDTH)),
    4681 => std_logic_vector(to_unsigned(6599, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4682 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4683 => std_logic_vector(to_unsigned(4597, LDPC_TABLE_DATA_WIDTH)),
    4684 => std_logic_vector(to_unsigned(4870, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4685 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4686 => std_logic_vector(to_unsigned(1228, LDPC_TABLE_DATA_WIDTH)),
    4687 => std_logic_vector(to_unsigned(6913, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4688 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4689 => std_logic_vector(to_unsigned(4159, LDPC_TABLE_DATA_WIDTH)),
    4690 => std_logic_vector(to_unsigned(1037, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4691 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4692 => std_logic_vector(to_unsigned(2916, LDPC_TABLE_DATA_WIDTH)),
    4693 => std_logic_vector(to_unsigned(2362, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4694 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4695 => std_logic_vector(to_unsigned(395, LDPC_TABLE_DATA_WIDTH)),
    4696 => std_logic_vector(to_unsigned(1226, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4697 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4698 => std_logic_vector(to_unsigned(6911, LDPC_TABLE_DATA_WIDTH)),
    4699 => std_logic_vector(to_unsigned(4548, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4700 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4701 => std_logic_vector(to_unsigned(4618, LDPC_TABLE_DATA_WIDTH)),
    4702 => std_logic_vector(to_unsigned(2241, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4703 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4704 => std_logic_vector(to_unsigned(4120, LDPC_TABLE_DATA_WIDTH)),
    4705 => std_logic_vector(to_unsigned(4280, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4706 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4707 => std_logic_vector(to_unsigned(5825, LDPC_TABLE_DATA_WIDTH)),
    4708 => std_logic_vector(to_unsigned(474, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4709 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4710 => std_logic_vector(to_unsigned(2154, LDPC_TABLE_DATA_WIDTH)),
    4711 => std_logic_vector(to_unsigned(5558, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4712 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4713 => std_logic_vector(to_unsigned(3793, LDPC_TABLE_DATA_WIDTH)),
    4714 => std_logic_vector(to_unsigned(5471, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4715 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4716 => std_logic_vector(to_unsigned(5707, LDPC_TABLE_DATA_WIDTH)),
    4717 => std_logic_vector(to_unsigned(1595, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4718 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4719 => std_logic_vector(to_unsigned(1403, LDPC_TABLE_DATA_WIDTH)),
    4720 => std_logic_vector(to_unsigned(325, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4721 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4722 => std_logic_vector(to_unsigned(6601, LDPC_TABLE_DATA_WIDTH)),
    4723 => std_logic_vector(to_unsigned(5183, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4724 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4725 => std_logic_vector(to_unsigned(6369, LDPC_TABLE_DATA_WIDTH)),
    4726 => std_logic_vector(to_unsigned(4569, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4727 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4728 => std_logic_vector(to_unsigned(4846, LDPC_TABLE_DATA_WIDTH)),
    4729 => std_logic_vector(to_unsigned(896, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4730 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4731 => std_logic_vector(to_unsigned(7092, LDPC_TABLE_DATA_WIDTH)),
    4732 => std_logic_vector(to_unsigned(6184, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4733 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4734 => std_logic_vector(to_unsigned(6764, LDPC_TABLE_DATA_WIDTH)),
    4735 => std_logic_vector(to_unsigned(7127, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4736 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4737 => std_logic_vector(to_unsigned(6358, LDPC_TABLE_DATA_WIDTH)),
    4738 => std_logic_vector(to_unsigned(1951, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4739 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4740 => std_logic_vector(to_unsigned(3117, LDPC_TABLE_DATA_WIDTH)),
    4741 => std_logic_vector(to_unsigned(6960, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4742 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4743 => std_logic_vector(to_unsigned(2710, LDPC_TABLE_DATA_WIDTH)),
    4744 => std_logic_vector(to_unsigned(7062, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4745 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4746 => std_logic_vector(to_unsigned(1133, LDPC_TABLE_DATA_WIDTH)),
    4747 => std_logic_vector(to_unsigned(3604, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4748 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4749 => std_logic_vector(to_unsigned(3694, LDPC_TABLE_DATA_WIDTH)),
    4750 => std_logic_vector(to_unsigned(657, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4751 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4752 => std_logic_vector(to_unsigned(1355, LDPC_TABLE_DATA_WIDTH)),
    4753 => std_logic_vector(to_unsigned(110, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4754 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4755 => std_logic_vector(to_unsigned(3329, LDPC_TABLE_DATA_WIDTH)),
    4756 => std_logic_vector(to_unsigned(6736, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4757 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4758 => std_logic_vector(to_unsigned(2505, LDPC_TABLE_DATA_WIDTH)),
    4759 => std_logic_vector(to_unsigned(3407, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4760 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4761 => std_logic_vector(to_unsigned(2462, LDPC_TABLE_DATA_WIDTH)),
    4762 => std_logic_vector(to_unsigned(4806, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4763 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4764 => std_logic_vector(to_unsigned(4216, LDPC_TABLE_DATA_WIDTH)),
    4765 => std_logic_vector(to_unsigned(214, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4766 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4767 => std_logic_vector(to_unsigned(5348, LDPC_TABLE_DATA_WIDTH)),
    4768 => std_logic_vector(to_unsigned(5619, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4769 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4770 => std_logic_vector(to_unsigned(6627, LDPC_TABLE_DATA_WIDTH)),
    4771 => std_logic_vector(to_unsigned(6243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4772 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4773 => std_logic_vector(to_unsigned(2644, LDPC_TABLE_DATA_WIDTH)),
    4774 => std_logic_vector(to_unsigned(5073, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4775 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4776 => std_logic_vector(to_unsigned(4212, LDPC_TABLE_DATA_WIDTH)),
    4777 => std_logic_vector(to_unsigned(5088, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4778 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4779 => std_logic_vector(to_unsigned(3463, LDPC_TABLE_DATA_WIDTH)),
    4780 => std_logic_vector(to_unsigned(3889, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4781 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4782 => std_logic_vector(to_unsigned(5306, LDPC_TABLE_DATA_WIDTH)),
    4783 => std_logic_vector(to_unsigned(478, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4784 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4785 => std_logic_vector(to_unsigned(4320, LDPC_TABLE_DATA_WIDTH)),
    4786 => std_logic_vector(to_unsigned(6121, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4787 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4788 => std_logic_vector(to_unsigned(3961, LDPC_TABLE_DATA_WIDTH)),
    4789 => std_logic_vector(to_unsigned(1125, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4790 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4791 => std_logic_vector(to_unsigned(5699, LDPC_TABLE_DATA_WIDTH)),
    4792 => std_logic_vector(to_unsigned(1195, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4793 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4794 => std_logic_vector(to_unsigned(6511, LDPC_TABLE_DATA_WIDTH)),
    4795 => std_logic_vector(to_unsigned(792, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4796 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4797 => std_logic_vector(to_unsigned(3934, LDPC_TABLE_DATA_WIDTH)),
    4798 => std_logic_vector(to_unsigned(2778, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4799 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4800 => std_logic_vector(to_unsigned(3238, LDPC_TABLE_DATA_WIDTH)),
    4801 => std_logic_vector(to_unsigned(6587, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4802 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4803 => std_logic_vector(to_unsigned(1111, LDPC_TABLE_DATA_WIDTH)),
    4804 => std_logic_vector(to_unsigned(6596, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4805 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4806 => std_logic_vector(to_unsigned(1457, LDPC_TABLE_DATA_WIDTH)),
    4807 => std_logic_vector(to_unsigned(6226, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4808 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4809 => std_logic_vector(to_unsigned(1446, LDPC_TABLE_DATA_WIDTH)),
    4810 => std_logic_vector(to_unsigned(3885, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4811 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4812 => std_logic_vector(to_unsigned(3907, LDPC_TABLE_DATA_WIDTH)),
    4813 => std_logic_vector(to_unsigned(4043, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4814 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4815 => std_logic_vector(to_unsigned(6839, LDPC_TABLE_DATA_WIDTH)),
    4816 => std_logic_vector(to_unsigned(2873, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4817 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4818 => std_logic_vector(to_unsigned(1733, LDPC_TABLE_DATA_WIDTH)),
    4819 => std_logic_vector(to_unsigned(5615, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4820 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4821 => std_logic_vector(to_unsigned(5202, LDPC_TABLE_DATA_WIDTH)),
    4822 => std_logic_vector(to_unsigned(4269, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4823 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4824 => std_logic_vector(to_unsigned(3024, LDPC_TABLE_DATA_WIDTH)),
    4825 => std_logic_vector(to_unsigned(4722, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4826 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4827 => std_logic_vector(to_unsigned(5445, LDPC_TABLE_DATA_WIDTH)),
    4828 => std_logic_vector(to_unsigned(6372, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4829 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4830 => std_logic_vector(to_unsigned(370, LDPC_TABLE_DATA_WIDTH)),
    4831 => std_logic_vector(to_unsigned(1828, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4832 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4833 => std_logic_vector(to_unsigned(4695, LDPC_TABLE_DATA_WIDTH)),
    4834 => std_logic_vector(to_unsigned(1600, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4835 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4836 => std_logic_vector(to_unsigned(680, LDPC_TABLE_DATA_WIDTH)),
    4837 => std_logic_vector(to_unsigned(2074, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4838 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4839 => std_logic_vector(to_unsigned(1801, LDPC_TABLE_DATA_WIDTH)),
    4840 => std_logic_vector(to_unsigned(6690, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4841 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4842 => std_logic_vector(to_unsigned(2669, LDPC_TABLE_DATA_WIDTH)),
    4843 => std_logic_vector(to_unsigned(1377, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4844 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4845 => std_logic_vector(to_unsigned(2463, LDPC_TABLE_DATA_WIDTH)),
    4846 => std_logic_vector(to_unsigned(1681, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4847 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4848 => std_logic_vector(to_unsigned(5972, LDPC_TABLE_DATA_WIDTH)),
    4849 => std_logic_vector(to_unsigned(5171, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4850 => std_logic_vector(to_unsigned(18, LDPC_TABLE_DATA_WIDTH)),
    4851 => std_logic_vector(to_unsigned(5728, LDPC_TABLE_DATA_WIDTH)),
    4852 => std_logic_vector(to_unsigned(4284, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4853 => std_logic_vector(to_unsigned(19, LDPC_TABLE_DATA_WIDTH)),
    4854 => std_logic_vector(to_unsigned(1696, LDPC_TABLE_DATA_WIDTH)),
    4855 => std_logic_vector(to_unsigned(1459, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_normal, C9_10
    4856 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4857 => std_logic_vector(to_unsigned(5611, LDPC_TABLE_DATA_WIDTH)),
    4858 => std_logic_vector(to_unsigned(2563, LDPC_TABLE_DATA_WIDTH)),
    4859 => std_logic_vector(to_unsigned(2900, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4860 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4861 => std_logic_vector(to_unsigned(5220, LDPC_TABLE_DATA_WIDTH)),
    4862 => std_logic_vector(to_unsigned(3143, LDPC_TABLE_DATA_WIDTH)),
    4863 => std_logic_vector(to_unsigned(4813, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4864 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4865 => std_logic_vector(to_unsigned(2481, LDPC_TABLE_DATA_WIDTH)),
    4866 => std_logic_vector(to_unsigned(834, LDPC_TABLE_DATA_WIDTH)),
    4867 => std_logic_vector(to_unsigned(81, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4868 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4869 => std_logic_vector(to_unsigned(6265, LDPC_TABLE_DATA_WIDTH)),
    4870 => std_logic_vector(to_unsigned(4064, LDPC_TABLE_DATA_WIDTH)),
    4871 => std_logic_vector(to_unsigned(4265, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4872 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4873 => std_logic_vector(to_unsigned(1055, LDPC_TABLE_DATA_WIDTH)),
    4874 => std_logic_vector(to_unsigned(2914, LDPC_TABLE_DATA_WIDTH)),
    4875 => std_logic_vector(to_unsigned(5638, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4876 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4877 => std_logic_vector(to_unsigned(1734, LDPC_TABLE_DATA_WIDTH)),
    4878 => std_logic_vector(to_unsigned(2182, LDPC_TABLE_DATA_WIDTH)),
    4879 => std_logic_vector(to_unsigned(3315, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4880 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4881 => std_logic_vector(to_unsigned(3342, LDPC_TABLE_DATA_WIDTH)),
    4882 => std_logic_vector(to_unsigned(5678, LDPC_TABLE_DATA_WIDTH)),
    4883 => std_logic_vector(to_unsigned(2246, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4884 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4885 => std_logic_vector(to_unsigned(2185, LDPC_TABLE_DATA_WIDTH)),
    4886 => std_logic_vector(to_unsigned(552, LDPC_TABLE_DATA_WIDTH)),
    4887 => std_logic_vector(to_unsigned(3385, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4888 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4889 => std_logic_vector(to_unsigned(2615, LDPC_TABLE_DATA_WIDTH)),
    4890 => std_logic_vector(to_unsigned(236, LDPC_TABLE_DATA_WIDTH)),
    4891 => std_logic_vector(to_unsigned(5334, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4892 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4893 => std_logic_vector(to_unsigned(1546, LDPC_TABLE_DATA_WIDTH)),
    4894 => std_logic_vector(to_unsigned(1755, LDPC_TABLE_DATA_WIDTH)),
    4895 => std_logic_vector(to_unsigned(3846, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4896 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4897 => std_logic_vector(to_unsigned(4154, LDPC_TABLE_DATA_WIDTH)),
    4898 => std_logic_vector(to_unsigned(5561, LDPC_TABLE_DATA_WIDTH)),
    4899 => std_logic_vector(to_unsigned(3142, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4900 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4901 => std_logic_vector(to_unsigned(4382, LDPC_TABLE_DATA_WIDTH)),
    4902 => std_logic_vector(to_unsigned(2957, LDPC_TABLE_DATA_WIDTH)),
    4903 => std_logic_vector(to_unsigned(5400, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4904 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4905 => std_logic_vector(to_unsigned(1209, LDPC_TABLE_DATA_WIDTH)),
    4906 => std_logic_vector(to_unsigned(5329, LDPC_TABLE_DATA_WIDTH)),
    4907 => std_logic_vector(to_unsigned(3179, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4908 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4909 => std_logic_vector(to_unsigned(1421, LDPC_TABLE_DATA_WIDTH)),
    4910 => std_logic_vector(to_unsigned(3528, LDPC_TABLE_DATA_WIDTH)),
    4911 => std_logic_vector(to_unsigned(6063, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4912 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4913 => std_logic_vector(to_unsigned(1480, LDPC_TABLE_DATA_WIDTH)),
    4914 => std_logic_vector(to_unsigned(1072, LDPC_TABLE_DATA_WIDTH)),
    4915 => std_logic_vector(to_unsigned(5398, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4916 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4917 => std_logic_vector(to_unsigned(3843, LDPC_TABLE_DATA_WIDTH)),
    4918 => std_logic_vector(to_unsigned(1777, LDPC_TABLE_DATA_WIDTH)),
    4919 => std_logic_vector(to_unsigned(4369, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4920 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4921 => std_logic_vector(to_unsigned(1334, LDPC_TABLE_DATA_WIDTH)),
    4922 => std_logic_vector(to_unsigned(2145, LDPC_TABLE_DATA_WIDTH)),
    4923 => std_logic_vector(to_unsigned(4163, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4924 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4925 => std_logic_vector(to_unsigned(2368, LDPC_TABLE_DATA_WIDTH)),
    4926 => std_logic_vector(to_unsigned(5055, LDPC_TABLE_DATA_WIDTH)),
    4927 => std_logic_vector(to_unsigned(260, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4928 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4929 => std_logic_vector(to_unsigned(6118, LDPC_TABLE_DATA_WIDTH)),
    4930 => std_logic_vector(to_unsigned(5405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4931 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4932 => std_logic_vector(to_unsigned(2994, LDPC_TABLE_DATA_WIDTH)),
    4933 => std_logic_vector(to_unsigned(4370, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4934 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4935 => std_logic_vector(to_unsigned(3405, LDPC_TABLE_DATA_WIDTH)),
    4936 => std_logic_vector(to_unsigned(1669, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4937 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4938 => std_logic_vector(to_unsigned(4640, LDPC_TABLE_DATA_WIDTH)),
    4939 => std_logic_vector(to_unsigned(5550, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4940 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4941 => std_logic_vector(to_unsigned(1354, LDPC_TABLE_DATA_WIDTH)),
    4942 => std_logic_vector(to_unsigned(3921, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4943 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4944 => std_logic_vector(to_unsigned(117, LDPC_TABLE_DATA_WIDTH)),
    4945 => std_logic_vector(to_unsigned(1713, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4946 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    4947 => std_logic_vector(to_unsigned(5425, LDPC_TABLE_DATA_WIDTH)),
    4948 => std_logic_vector(to_unsigned(2866, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4949 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    4950 => std_logic_vector(to_unsigned(6047, LDPC_TABLE_DATA_WIDTH)),
    4951 => std_logic_vector(to_unsigned(683, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4952 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    4953 => std_logic_vector(to_unsigned(5616, LDPC_TABLE_DATA_WIDTH)),
    4954 => std_logic_vector(to_unsigned(2582, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4955 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    4956 => std_logic_vector(to_unsigned(2108, LDPC_TABLE_DATA_WIDTH)),
    4957 => std_logic_vector(to_unsigned(1179, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4958 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    4959 => std_logic_vector(to_unsigned(933, LDPC_TABLE_DATA_WIDTH)),
    4960 => std_logic_vector(to_unsigned(4921, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4961 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    4962 => std_logic_vector(to_unsigned(5953, LDPC_TABLE_DATA_WIDTH)),
    4963 => std_logic_vector(to_unsigned(2261, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4964 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    4965 => std_logic_vector(to_unsigned(1430, LDPC_TABLE_DATA_WIDTH)),
    4966 => std_logic_vector(to_unsigned(4699, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4967 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    4968 => std_logic_vector(to_unsigned(5905, LDPC_TABLE_DATA_WIDTH)),
    4969 => std_logic_vector(to_unsigned(480, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4970 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    4971 => std_logic_vector(to_unsigned(4289, LDPC_TABLE_DATA_WIDTH)),
    4972 => std_logic_vector(to_unsigned(1846, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4973 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    4974 => std_logic_vector(to_unsigned(5374, LDPC_TABLE_DATA_WIDTH)),
    4975 => std_logic_vector(to_unsigned(6208, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4976 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    4977 => std_logic_vector(to_unsigned(1775, LDPC_TABLE_DATA_WIDTH)),
    4978 => std_logic_vector(to_unsigned(3476, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4979 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    4980 => std_logic_vector(to_unsigned(3216, LDPC_TABLE_DATA_WIDTH)),
    4981 => std_logic_vector(to_unsigned(2178, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4982 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    4983 => std_logic_vector(to_unsigned(4165, LDPC_TABLE_DATA_WIDTH)),
    4984 => std_logic_vector(to_unsigned(884, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4985 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    4986 => std_logic_vector(to_unsigned(2896, LDPC_TABLE_DATA_WIDTH)),
    4987 => std_logic_vector(to_unsigned(3744, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4988 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    4989 => std_logic_vector(to_unsigned(874, LDPC_TABLE_DATA_WIDTH)),
    4990 => std_logic_vector(to_unsigned(2801, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4991 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    4992 => std_logic_vector(to_unsigned(3423, LDPC_TABLE_DATA_WIDTH)),
    4993 => std_logic_vector(to_unsigned(5579, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4994 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    4995 => std_logic_vector(to_unsigned(3404, LDPC_TABLE_DATA_WIDTH)),
    4996 => std_logic_vector(to_unsigned(3552, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    4997 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    4998 => std_logic_vector(to_unsigned(2876, LDPC_TABLE_DATA_WIDTH)),
    4999 => std_logic_vector(to_unsigned(5515, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5000 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5001 => std_logic_vector(to_unsigned(516, LDPC_TABLE_DATA_WIDTH)),
    5002 => std_logic_vector(to_unsigned(1719, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5003 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5004 => std_logic_vector(to_unsigned(765, LDPC_TABLE_DATA_WIDTH)),
    5005 => std_logic_vector(to_unsigned(3631, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5006 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5007 => std_logic_vector(to_unsigned(5059, LDPC_TABLE_DATA_WIDTH)),
    5008 => std_logic_vector(to_unsigned(1441, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5009 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5010 => std_logic_vector(to_unsigned(5629, LDPC_TABLE_DATA_WIDTH)),
    5011 => std_logic_vector(to_unsigned(598, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5012 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5013 => std_logic_vector(to_unsigned(5405, LDPC_TABLE_DATA_WIDTH)),
    5014 => std_logic_vector(to_unsigned(473, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5015 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5016 => std_logic_vector(to_unsigned(4724, LDPC_TABLE_DATA_WIDTH)),
    5017 => std_logic_vector(to_unsigned(5210, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5018 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5019 => std_logic_vector(to_unsigned(155, LDPC_TABLE_DATA_WIDTH)),
    5020 => std_logic_vector(to_unsigned(1832, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5021 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5022 => std_logic_vector(to_unsigned(1689, LDPC_TABLE_DATA_WIDTH)),
    5023 => std_logic_vector(to_unsigned(2229, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5024 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5025 => std_logic_vector(to_unsigned(449, LDPC_TABLE_DATA_WIDTH)),
    5026 => std_logic_vector(to_unsigned(1164, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5027 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5028 => std_logic_vector(to_unsigned(2308, LDPC_TABLE_DATA_WIDTH)),
    5029 => std_logic_vector(to_unsigned(3088, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5030 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5031 => std_logic_vector(to_unsigned(1122, LDPC_TABLE_DATA_WIDTH)),
    5032 => std_logic_vector(to_unsigned(669, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5033 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5034 => std_logic_vector(to_unsigned(2268, LDPC_TABLE_DATA_WIDTH)),
    5035 => std_logic_vector(to_unsigned(5758, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5036 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5037 => std_logic_vector(to_unsigned(5878, LDPC_TABLE_DATA_WIDTH)),
    5038 => std_logic_vector(to_unsigned(2609, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5039 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5040 => std_logic_vector(to_unsigned(782, LDPC_TABLE_DATA_WIDTH)),
    5041 => std_logic_vector(to_unsigned(3359, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5042 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5043 => std_logic_vector(to_unsigned(1231, LDPC_TABLE_DATA_WIDTH)),
    5044 => std_logic_vector(to_unsigned(4231, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5045 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5046 => std_logic_vector(to_unsigned(4225, LDPC_TABLE_DATA_WIDTH)),
    5047 => std_logic_vector(to_unsigned(2052, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5048 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5049 => std_logic_vector(to_unsigned(4286, LDPC_TABLE_DATA_WIDTH)),
    5050 => std_logic_vector(to_unsigned(3517, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5051 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5052 => std_logic_vector(to_unsigned(5531, LDPC_TABLE_DATA_WIDTH)),
    5053 => std_logic_vector(to_unsigned(3184, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5054 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5055 => std_logic_vector(to_unsigned(1935, LDPC_TABLE_DATA_WIDTH)),
    5056 => std_logic_vector(to_unsigned(4560, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5057 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5058 => std_logic_vector(to_unsigned(1174, LDPC_TABLE_DATA_WIDTH)),
    5059 => std_logic_vector(to_unsigned(131, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5060 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5061 => std_logic_vector(to_unsigned(3115, LDPC_TABLE_DATA_WIDTH)),
    5062 => std_logic_vector(to_unsigned(956, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5063 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5064 => std_logic_vector(to_unsigned(3129, LDPC_TABLE_DATA_WIDTH)),
    5065 => std_logic_vector(to_unsigned(1088, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5066 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5067 => std_logic_vector(to_unsigned(5238, LDPC_TABLE_DATA_WIDTH)),
    5068 => std_logic_vector(to_unsigned(4440, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5069 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5070 => std_logic_vector(to_unsigned(5722, LDPC_TABLE_DATA_WIDTH)),
    5071 => std_logic_vector(to_unsigned(4280, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5072 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5073 => std_logic_vector(to_unsigned(3540, LDPC_TABLE_DATA_WIDTH)),
    5074 => std_logic_vector(to_unsigned(375, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5075 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5076 => std_logic_vector(to_unsigned(191, LDPC_TABLE_DATA_WIDTH)),
    5077 => std_logic_vector(to_unsigned(2782, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5078 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5079 => std_logic_vector(to_unsigned(906, LDPC_TABLE_DATA_WIDTH)),
    5080 => std_logic_vector(to_unsigned(4432, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5081 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5082 => std_logic_vector(to_unsigned(3225, LDPC_TABLE_DATA_WIDTH)),
    5083 => std_logic_vector(to_unsigned(1111, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5084 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5085 => std_logic_vector(to_unsigned(6296, LDPC_TABLE_DATA_WIDTH)),
    5086 => std_logic_vector(to_unsigned(2583, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5087 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5088 => std_logic_vector(to_unsigned(1457, LDPC_TABLE_DATA_WIDTH)),
    5089 => std_logic_vector(to_unsigned(903, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5090 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5091 => std_logic_vector(to_unsigned(855, LDPC_TABLE_DATA_WIDTH)),
    5092 => std_logic_vector(to_unsigned(4475, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5093 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5094 => std_logic_vector(to_unsigned(4097, LDPC_TABLE_DATA_WIDTH)),
    5095 => std_logic_vector(to_unsigned(3970, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5096 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5097 => std_logic_vector(to_unsigned(4433, LDPC_TABLE_DATA_WIDTH)),
    5098 => std_logic_vector(to_unsigned(4361, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5099 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5100 => std_logic_vector(to_unsigned(5198, LDPC_TABLE_DATA_WIDTH)),
    5101 => std_logic_vector(to_unsigned(541, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5102 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5103 => std_logic_vector(to_unsigned(1146, LDPC_TABLE_DATA_WIDTH)),
    5104 => std_logic_vector(to_unsigned(4426, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5105 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5106 => std_logic_vector(to_unsigned(3202, LDPC_TABLE_DATA_WIDTH)),
    5107 => std_logic_vector(to_unsigned(2902, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5108 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5109 => std_logic_vector(to_unsigned(2724, LDPC_TABLE_DATA_WIDTH)),
    5110 => std_logic_vector(to_unsigned(525, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5111 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5112 => std_logic_vector(to_unsigned(1083, LDPC_TABLE_DATA_WIDTH)),
    5113 => std_logic_vector(to_unsigned(4124, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5114 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5115 => std_logic_vector(to_unsigned(2326, LDPC_TABLE_DATA_WIDTH)),
    5116 => std_logic_vector(to_unsigned(6003, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5117 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5118 => std_logic_vector(to_unsigned(5605, LDPC_TABLE_DATA_WIDTH)),
    5119 => std_logic_vector(to_unsigned(5990, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5120 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5121 => std_logic_vector(to_unsigned(4376, LDPC_TABLE_DATA_WIDTH)),
    5122 => std_logic_vector(to_unsigned(1579, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5123 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5124 => std_logic_vector(to_unsigned(4407, LDPC_TABLE_DATA_WIDTH)),
    5125 => std_logic_vector(to_unsigned(984, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5126 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5127 => std_logic_vector(to_unsigned(1332, LDPC_TABLE_DATA_WIDTH)),
    5128 => std_logic_vector(to_unsigned(6163, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5129 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5130 => std_logic_vector(to_unsigned(5359, LDPC_TABLE_DATA_WIDTH)),
    5131 => std_logic_vector(to_unsigned(3975, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5132 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5133 => std_logic_vector(to_unsigned(1907, LDPC_TABLE_DATA_WIDTH)),
    5134 => std_logic_vector(to_unsigned(1854, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5135 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5136 => std_logic_vector(to_unsigned(3601, LDPC_TABLE_DATA_WIDTH)),
    5137 => std_logic_vector(to_unsigned(5748, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5138 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5139 => std_logic_vector(to_unsigned(6056, LDPC_TABLE_DATA_WIDTH)),
    5140 => std_logic_vector(to_unsigned(3266, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5141 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5142 => std_logic_vector(to_unsigned(3322, LDPC_TABLE_DATA_WIDTH)),
    5143 => std_logic_vector(to_unsigned(4085, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5144 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5145 => std_logic_vector(to_unsigned(1768, LDPC_TABLE_DATA_WIDTH)),
    5146 => std_logic_vector(to_unsigned(3244, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5147 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5148 => std_logic_vector(to_unsigned(2149, LDPC_TABLE_DATA_WIDTH)),
    5149 => std_logic_vector(to_unsigned(144, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5150 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5151 => std_logic_vector(to_unsigned(1589, LDPC_TABLE_DATA_WIDTH)),
    5152 => std_logic_vector(to_unsigned(4291, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5153 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5154 => std_logic_vector(to_unsigned(5154, LDPC_TABLE_DATA_WIDTH)),
    5155 => std_logic_vector(to_unsigned(1252, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5156 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5157 => std_logic_vector(to_unsigned(1855, LDPC_TABLE_DATA_WIDTH)),
    5158 => std_logic_vector(to_unsigned(5939, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5159 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5160 => std_logic_vector(to_unsigned(4820, LDPC_TABLE_DATA_WIDTH)),
    5161 => std_logic_vector(to_unsigned(2706, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5162 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5163 => std_logic_vector(to_unsigned(1475, LDPC_TABLE_DATA_WIDTH)),
    5164 => std_logic_vector(to_unsigned(3360, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5165 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5166 => std_logic_vector(to_unsigned(4266, LDPC_TABLE_DATA_WIDTH)),
    5167 => std_logic_vector(to_unsigned(693, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5168 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5169 => std_logic_vector(to_unsigned(4156, LDPC_TABLE_DATA_WIDTH)),
    5170 => std_logic_vector(to_unsigned(2018, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5171 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5172 => std_logic_vector(to_unsigned(2103, LDPC_TABLE_DATA_WIDTH)),
    5173 => std_logic_vector(to_unsigned(752, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5174 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5175 => std_logic_vector(to_unsigned(3710, LDPC_TABLE_DATA_WIDTH)),
    5176 => std_logic_vector(to_unsigned(3853, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5177 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5178 => std_logic_vector(to_unsigned(5123, LDPC_TABLE_DATA_WIDTH)),
    5179 => std_logic_vector(to_unsigned(931, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5180 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5181 => std_logic_vector(to_unsigned(6146, LDPC_TABLE_DATA_WIDTH)),
    5182 => std_logic_vector(to_unsigned(3323, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5183 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5184 => std_logic_vector(to_unsigned(1939, LDPC_TABLE_DATA_WIDTH)),
    5185 => std_logic_vector(to_unsigned(5002, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5186 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5187 => std_logic_vector(to_unsigned(5140, LDPC_TABLE_DATA_WIDTH)),
    5188 => std_logic_vector(to_unsigned(1437, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5189 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5190 => std_logic_vector(to_unsigned(1263, LDPC_TABLE_DATA_WIDTH)),
    5191 => std_logic_vector(to_unsigned(293, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5192 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5193 => std_logic_vector(to_unsigned(5949, LDPC_TABLE_DATA_WIDTH)),
    5194 => std_logic_vector(to_unsigned(4665, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5195 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5196 => std_logic_vector(to_unsigned(4548, LDPC_TABLE_DATA_WIDTH)),
    5197 => std_logic_vector(to_unsigned(6380, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5198 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5199 => std_logic_vector(to_unsigned(3171, LDPC_TABLE_DATA_WIDTH)),
    5200 => std_logic_vector(to_unsigned(4690, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5201 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5202 => std_logic_vector(to_unsigned(5204, LDPC_TABLE_DATA_WIDTH)),
    5203 => std_logic_vector(to_unsigned(2114, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5204 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5205 => std_logic_vector(to_unsigned(6384, LDPC_TABLE_DATA_WIDTH)),
    5206 => std_logic_vector(to_unsigned(5565, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5207 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5208 => std_logic_vector(to_unsigned(5722, LDPC_TABLE_DATA_WIDTH)),
    5209 => std_logic_vector(to_unsigned(1757, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5210 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5211 => std_logic_vector(to_unsigned(2805, LDPC_TABLE_DATA_WIDTH)),
    5212 => std_logic_vector(to_unsigned(6264, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5213 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5214 => std_logic_vector(to_unsigned(1202, LDPC_TABLE_DATA_WIDTH)),
    5215 => std_logic_vector(to_unsigned(2616, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5216 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5217 => std_logic_vector(to_unsigned(1018, LDPC_TABLE_DATA_WIDTH)),
    5218 => std_logic_vector(to_unsigned(3244, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5219 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5220 => std_logic_vector(to_unsigned(4018, LDPC_TABLE_DATA_WIDTH)),
    5221 => std_logic_vector(to_unsigned(5289, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5222 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5223 => std_logic_vector(to_unsigned(2257, LDPC_TABLE_DATA_WIDTH)),
    5224 => std_logic_vector(to_unsigned(3067, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5225 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5226 => std_logic_vector(to_unsigned(2483, LDPC_TABLE_DATA_WIDTH)),
    5227 => std_logic_vector(to_unsigned(3073, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5228 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5229 => std_logic_vector(to_unsigned(1196, LDPC_TABLE_DATA_WIDTH)),
    5230 => std_logic_vector(to_unsigned(5329, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5231 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5232 => std_logic_vector(to_unsigned(649, LDPC_TABLE_DATA_WIDTH)),
    5233 => std_logic_vector(to_unsigned(3918, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5234 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5235 => std_logic_vector(to_unsigned(3791, LDPC_TABLE_DATA_WIDTH)),
    5236 => std_logic_vector(to_unsigned(4581, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5237 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5238 => std_logic_vector(to_unsigned(5028, LDPC_TABLE_DATA_WIDTH)),
    5239 => std_logic_vector(to_unsigned(3803, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5240 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5241 => std_logic_vector(to_unsigned(3119, LDPC_TABLE_DATA_WIDTH)),
    5242 => std_logic_vector(to_unsigned(3506, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5243 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5244 => std_logic_vector(to_unsigned(4779, LDPC_TABLE_DATA_WIDTH)),
    5245 => std_logic_vector(to_unsigned(431, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5246 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5247 => std_logic_vector(to_unsigned(3888, LDPC_TABLE_DATA_WIDTH)),
    5248 => std_logic_vector(to_unsigned(5510, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5249 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5250 => std_logic_vector(to_unsigned(4387, LDPC_TABLE_DATA_WIDTH)),
    5251 => std_logic_vector(to_unsigned(4084, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5252 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5253 => std_logic_vector(to_unsigned(5836, LDPC_TABLE_DATA_WIDTH)),
    5254 => std_logic_vector(to_unsigned(1692, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5255 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5256 => std_logic_vector(to_unsigned(5126, LDPC_TABLE_DATA_WIDTH)),
    5257 => std_logic_vector(to_unsigned(1078, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5258 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5259 => std_logic_vector(to_unsigned(5721, LDPC_TABLE_DATA_WIDTH)),
    5260 => std_logic_vector(to_unsigned(6165, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5261 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5262 => std_logic_vector(to_unsigned(3540, LDPC_TABLE_DATA_WIDTH)),
    5263 => std_logic_vector(to_unsigned(2499, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5264 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5265 => std_logic_vector(to_unsigned(2225, LDPC_TABLE_DATA_WIDTH)),
    5266 => std_logic_vector(to_unsigned(6348, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5267 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5268 => std_logic_vector(to_unsigned(1044, LDPC_TABLE_DATA_WIDTH)),
    5269 => std_logic_vector(to_unsigned(1484, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5270 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5271 => std_logic_vector(to_unsigned(6323, LDPC_TABLE_DATA_WIDTH)),
    5272 => std_logic_vector(to_unsigned(4042, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5273 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5274 => std_logic_vector(to_unsigned(1313, LDPC_TABLE_DATA_WIDTH)),
    5275 => std_logic_vector(to_unsigned(5603, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5276 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5277 => std_logic_vector(to_unsigned(1303, LDPC_TABLE_DATA_WIDTH)),
    5278 => std_logic_vector(to_unsigned(3496, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5279 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5280 => std_logic_vector(to_unsigned(3516, LDPC_TABLE_DATA_WIDTH)),
    5281 => std_logic_vector(to_unsigned(3639, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5282 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5283 => std_logic_vector(to_unsigned(5161, LDPC_TABLE_DATA_WIDTH)),
    5284 => std_logic_vector(to_unsigned(2293, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5285 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5286 => std_logic_vector(to_unsigned(4682, LDPC_TABLE_DATA_WIDTH)),
    5287 => std_logic_vector(to_unsigned(3845, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5288 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5289 => std_logic_vector(to_unsigned(3045, LDPC_TABLE_DATA_WIDTH)),
    5290 => std_logic_vector(to_unsigned(643, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5291 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5292 => std_logic_vector(to_unsigned(2818, LDPC_TABLE_DATA_WIDTH)),
    5293 => std_logic_vector(to_unsigned(2616, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5294 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5295 => std_logic_vector(to_unsigned(3267, LDPC_TABLE_DATA_WIDTH)),
    5296 => std_logic_vector(to_unsigned(649, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5297 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5298 => std_logic_vector(to_unsigned(6236, LDPC_TABLE_DATA_WIDTH)),
    5299 => std_logic_vector(to_unsigned(593, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5300 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5301 => std_logic_vector(to_unsigned(646, LDPC_TABLE_DATA_WIDTH)),
    5302 => std_logic_vector(to_unsigned(2948, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5303 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5304 => std_logic_vector(to_unsigned(4213, LDPC_TABLE_DATA_WIDTH)),
    5305 => std_logic_vector(to_unsigned(1442, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5306 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5307 => std_logic_vector(to_unsigned(5779, LDPC_TABLE_DATA_WIDTH)),
    5308 => std_logic_vector(to_unsigned(1596, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5309 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5310 => std_logic_vector(to_unsigned(2403, LDPC_TABLE_DATA_WIDTH)),
    5311 => std_logic_vector(to_unsigned(1237, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5312 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5313 => std_logic_vector(to_unsigned(2217, LDPC_TABLE_DATA_WIDTH)),
    5314 => std_logic_vector(to_unsigned(1514, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5315 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5316 => std_logic_vector(to_unsigned(5609, LDPC_TABLE_DATA_WIDTH)),
    5317 => std_logic_vector(to_unsigned(716, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5318 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5319 => std_logic_vector(to_unsigned(5155, LDPC_TABLE_DATA_WIDTH)),
    5320 => std_logic_vector(to_unsigned(3858, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5321 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5322 => std_logic_vector(to_unsigned(1517, LDPC_TABLE_DATA_WIDTH)),
    5323 => std_logic_vector(to_unsigned(1312, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5324 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5325 => std_logic_vector(to_unsigned(2554, LDPC_TABLE_DATA_WIDTH)),
    5326 => std_logic_vector(to_unsigned(3158, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5327 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5328 => std_logic_vector(to_unsigned(5280, LDPC_TABLE_DATA_WIDTH)),
    5329 => std_logic_vector(to_unsigned(2643, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5330 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5331 => std_logic_vector(to_unsigned(4990, LDPC_TABLE_DATA_WIDTH)),
    5332 => std_logic_vector(to_unsigned(1353, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5333 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5334 => std_logic_vector(to_unsigned(5648, LDPC_TABLE_DATA_WIDTH)),
    5335 => std_logic_vector(to_unsigned(1170, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5336 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5337 => std_logic_vector(to_unsigned(1152, LDPC_TABLE_DATA_WIDTH)),
    5338 => std_logic_vector(to_unsigned(4366, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5339 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5340 => std_logic_vector(to_unsigned(3561, LDPC_TABLE_DATA_WIDTH)),
    5341 => std_logic_vector(to_unsigned(5368, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5342 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5343 => std_logic_vector(to_unsigned(3581, LDPC_TABLE_DATA_WIDTH)),
    5344 => std_logic_vector(to_unsigned(1411, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5345 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5346 => std_logic_vector(to_unsigned(5647, LDPC_TABLE_DATA_WIDTH)),
    5347 => std_logic_vector(to_unsigned(4661, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5348 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5349 => std_logic_vector(to_unsigned(1542, LDPC_TABLE_DATA_WIDTH)),
    5350 => std_logic_vector(to_unsigned(5401, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5351 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    5352 => std_logic_vector(to_unsigned(5078, LDPC_TABLE_DATA_WIDTH)),
    5353 => std_logic_vector(to_unsigned(2687, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5354 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    5355 => std_logic_vector(to_unsigned(316, LDPC_TABLE_DATA_WIDTH)),
    5356 => std_logic_vector(to_unsigned(1755, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5357 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    5358 => std_logic_vector(to_unsigned(3392, LDPC_TABLE_DATA_WIDTH)),
    5359 => std_logic_vector(to_unsigned(1991, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C1_2
    5360 => std_logic_vector(to_unsigned(20, LDPC_TABLE_DATA_WIDTH)),
    5361 => std_logic_vector(to_unsigned(712, LDPC_TABLE_DATA_WIDTH)),
    5362 => std_logic_vector(to_unsigned(2386, LDPC_TABLE_DATA_WIDTH)),
    5363 => std_logic_vector(to_unsigned(6354, LDPC_TABLE_DATA_WIDTH)),
    5364 => std_logic_vector(to_unsigned(4061, LDPC_TABLE_DATA_WIDTH)),
    5365 => std_logic_vector(to_unsigned(1062, LDPC_TABLE_DATA_WIDTH)),
    5366 => std_logic_vector(to_unsigned(5045, LDPC_TABLE_DATA_WIDTH)),
    5367 => std_logic_vector(to_unsigned(5158, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5368 => std_logic_vector(to_unsigned(21, LDPC_TABLE_DATA_WIDTH)),
    5369 => std_logic_vector(to_unsigned(2543, LDPC_TABLE_DATA_WIDTH)),
    5370 => std_logic_vector(to_unsigned(5748, LDPC_TABLE_DATA_WIDTH)),
    5371 => std_logic_vector(to_unsigned(4822, LDPC_TABLE_DATA_WIDTH)),
    5372 => std_logic_vector(to_unsigned(2348, LDPC_TABLE_DATA_WIDTH)),
    5373 => std_logic_vector(to_unsigned(3089, LDPC_TABLE_DATA_WIDTH)),
    5374 => std_logic_vector(to_unsigned(6328, LDPC_TABLE_DATA_WIDTH)),
    5375 => std_logic_vector(to_unsigned(5876, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5376 => std_logic_vector(to_unsigned(22, LDPC_TABLE_DATA_WIDTH)),
    5377 => std_logic_vector(to_unsigned(926, LDPC_TABLE_DATA_WIDTH)),
    5378 => std_logic_vector(to_unsigned(5701, LDPC_TABLE_DATA_WIDTH)),
    5379 => std_logic_vector(to_unsigned(269, LDPC_TABLE_DATA_WIDTH)),
    5380 => std_logic_vector(to_unsigned(3693, LDPC_TABLE_DATA_WIDTH)),
    5381 => std_logic_vector(to_unsigned(2438, LDPC_TABLE_DATA_WIDTH)),
    5382 => std_logic_vector(to_unsigned(3190, LDPC_TABLE_DATA_WIDTH)),
    5383 => std_logic_vector(to_unsigned(3507, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5384 => std_logic_vector(to_unsigned(23, LDPC_TABLE_DATA_WIDTH)),
    5385 => std_logic_vector(to_unsigned(2802, LDPC_TABLE_DATA_WIDTH)),
    5386 => std_logic_vector(to_unsigned(4520, LDPC_TABLE_DATA_WIDTH)),
    5387 => std_logic_vector(to_unsigned(3577, LDPC_TABLE_DATA_WIDTH)),
    5388 => std_logic_vector(to_unsigned(5324, LDPC_TABLE_DATA_WIDTH)),
    5389 => std_logic_vector(to_unsigned(1091, LDPC_TABLE_DATA_WIDTH)),
    5390 => std_logic_vector(to_unsigned(4667, LDPC_TABLE_DATA_WIDTH)),
    5391 => std_logic_vector(to_unsigned(4449, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5392 => std_logic_vector(to_unsigned(24, LDPC_TABLE_DATA_WIDTH)),
    5393 => std_logic_vector(to_unsigned(5140, LDPC_TABLE_DATA_WIDTH)),
    5394 => std_logic_vector(to_unsigned(2003, LDPC_TABLE_DATA_WIDTH)),
    5395 => std_logic_vector(to_unsigned(1263, LDPC_TABLE_DATA_WIDTH)),
    5396 => std_logic_vector(to_unsigned(4742, LDPC_TABLE_DATA_WIDTH)),
    5397 => std_logic_vector(to_unsigned(6497, LDPC_TABLE_DATA_WIDTH)),
    5398 => std_logic_vector(to_unsigned(1185, LDPC_TABLE_DATA_WIDTH)),
    5399 => std_logic_vector(to_unsigned(6202, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5400 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5401 => std_logic_vector(to_unsigned(4046, LDPC_TABLE_DATA_WIDTH)),
    5402 => std_logic_vector(to_unsigned(6934, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5403 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5404 => std_logic_vector(to_unsigned(2855, LDPC_TABLE_DATA_WIDTH)),
    5405 => std_logic_vector(to_unsigned(66, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5406 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5407 => std_logic_vector(to_unsigned(6694, LDPC_TABLE_DATA_WIDTH)),
    5408 => std_logic_vector(to_unsigned(212, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5409 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5410 => std_logic_vector(to_unsigned(3439, LDPC_TABLE_DATA_WIDTH)),
    5411 => std_logic_vector(to_unsigned(1158, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5412 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5413 => std_logic_vector(to_unsigned(3850, LDPC_TABLE_DATA_WIDTH)),
    5414 => std_logic_vector(to_unsigned(4422, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5415 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5416 => std_logic_vector(to_unsigned(5924, LDPC_TABLE_DATA_WIDTH)),
    5417 => std_logic_vector(to_unsigned(290, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5418 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5419 => std_logic_vector(to_unsigned(1467, LDPC_TABLE_DATA_WIDTH)),
    5420 => std_logic_vector(to_unsigned(4049, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5421 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5422 => std_logic_vector(to_unsigned(7820, LDPC_TABLE_DATA_WIDTH)),
    5423 => std_logic_vector(to_unsigned(2242, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5424 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5425 => std_logic_vector(to_unsigned(4606, LDPC_TABLE_DATA_WIDTH)),
    5426 => std_logic_vector(to_unsigned(3080, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5427 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5428 => std_logic_vector(to_unsigned(4633, LDPC_TABLE_DATA_WIDTH)),
    5429 => std_logic_vector(to_unsigned(7877, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5430 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5431 => std_logic_vector(to_unsigned(3884, LDPC_TABLE_DATA_WIDTH)),
    5432 => std_logic_vector(to_unsigned(6868, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5433 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5434 => std_logic_vector(to_unsigned(8935, LDPC_TABLE_DATA_WIDTH)),
    5435 => std_logic_vector(to_unsigned(4996, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5436 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5437 => std_logic_vector(to_unsigned(3028, LDPC_TABLE_DATA_WIDTH)),
    5438 => std_logic_vector(to_unsigned(764, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5439 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5440 => std_logic_vector(to_unsigned(5988, LDPC_TABLE_DATA_WIDTH)),
    5441 => std_logic_vector(to_unsigned(1057, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5442 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5443 => std_logic_vector(to_unsigned(7411, LDPC_TABLE_DATA_WIDTH)),
    5444 => std_logic_vector(to_unsigned(3450, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C1_3
    5445 => std_logic_vector(to_unsigned(416, LDPC_TABLE_DATA_WIDTH)),
    5446 => std_logic_vector(to_unsigned(8909, LDPC_TABLE_DATA_WIDTH)),
    5447 => std_logic_vector(to_unsigned(4156, LDPC_TABLE_DATA_WIDTH)),
    5448 => std_logic_vector(to_unsigned(3216, LDPC_TABLE_DATA_WIDTH)),
    5449 => std_logic_vector(to_unsigned(3112, LDPC_TABLE_DATA_WIDTH)),
    5450 => std_logic_vector(to_unsigned(2560, LDPC_TABLE_DATA_WIDTH)),
    5451 => std_logic_vector(to_unsigned(2912, LDPC_TABLE_DATA_WIDTH)),
    5452 => std_logic_vector(to_unsigned(6405, LDPC_TABLE_DATA_WIDTH)),
    5453 => std_logic_vector(to_unsigned(8593, LDPC_TABLE_DATA_WIDTH)),
    5454 => std_logic_vector(to_unsigned(4969, LDPC_TABLE_DATA_WIDTH)),
    5455 => std_logic_vector(to_unsigned(6723, LDPC_TABLE_DATA_WIDTH)),
    5456 => std_logic_vector(to_unsigned(6912, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5457 => std_logic_vector(to_unsigned(8978, LDPC_TABLE_DATA_WIDTH)),
    5458 => std_logic_vector(to_unsigned(3011, LDPC_TABLE_DATA_WIDTH)),
    5459 => std_logic_vector(to_unsigned(4339, LDPC_TABLE_DATA_WIDTH)),
    5460 => std_logic_vector(to_unsigned(9312, LDPC_TABLE_DATA_WIDTH)),
    5461 => std_logic_vector(to_unsigned(6396, LDPC_TABLE_DATA_WIDTH)),
    5462 => std_logic_vector(to_unsigned(2957, LDPC_TABLE_DATA_WIDTH)),
    5463 => std_logic_vector(to_unsigned(7288, LDPC_TABLE_DATA_WIDTH)),
    5464 => std_logic_vector(to_unsigned(5485, LDPC_TABLE_DATA_WIDTH)),
    5465 => std_logic_vector(to_unsigned(6031, LDPC_TABLE_DATA_WIDTH)),
    5466 => std_logic_vector(to_unsigned(10218, LDPC_TABLE_DATA_WIDTH)),
    5467 => std_logic_vector(to_unsigned(2226, LDPC_TABLE_DATA_WIDTH)),
    5468 => std_logic_vector(to_unsigned(3575, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5469 => std_logic_vector(to_unsigned(3383, LDPC_TABLE_DATA_WIDTH)),
    5470 => std_logic_vector(to_unsigned(10059, LDPC_TABLE_DATA_WIDTH)),
    5471 => std_logic_vector(to_unsigned(1114, LDPC_TABLE_DATA_WIDTH)),
    5472 => std_logic_vector(to_unsigned(10008, LDPC_TABLE_DATA_WIDTH)),
    5473 => std_logic_vector(to_unsigned(10147, LDPC_TABLE_DATA_WIDTH)),
    5474 => std_logic_vector(to_unsigned(9384, LDPC_TABLE_DATA_WIDTH)),
    5475 => std_logic_vector(to_unsigned(4290, LDPC_TABLE_DATA_WIDTH)),
    5476 => std_logic_vector(to_unsigned(434, LDPC_TABLE_DATA_WIDTH)),
    5477 => std_logic_vector(to_unsigned(5139, LDPC_TABLE_DATA_WIDTH)),
    5478 => std_logic_vector(to_unsigned(3536, LDPC_TABLE_DATA_WIDTH)),
    5479 => std_logic_vector(to_unsigned(1965, LDPC_TABLE_DATA_WIDTH)),
    5480 => std_logic_vector(to_unsigned(2291, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5481 => std_logic_vector(to_unsigned(2797, LDPC_TABLE_DATA_WIDTH)),
    5482 => std_logic_vector(to_unsigned(3693, LDPC_TABLE_DATA_WIDTH)),
    5483 => std_logic_vector(to_unsigned(7615, LDPC_TABLE_DATA_WIDTH)),
    5484 => std_logic_vector(to_unsigned(7077, LDPC_TABLE_DATA_WIDTH)),
    5485 => std_logic_vector(to_unsigned(743, LDPC_TABLE_DATA_WIDTH)),
    5486 => std_logic_vector(to_unsigned(1941, LDPC_TABLE_DATA_WIDTH)),
    5487 => std_logic_vector(to_unsigned(8716, LDPC_TABLE_DATA_WIDTH)),
    5488 => std_logic_vector(to_unsigned(6215, LDPC_TABLE_DATA_WIDTH)),
    5489 => std_logic_vector(to_unsigned(3840, LDPC_TABLE_DATA_WIDTH)),
    5490 => std_logic_vector(to_unsigned(5140, LDPC_TABLE_DATA_WIDTH)),
    5491 => std_logic_vector(to_unsigned(4582, LDPC_TABLE_DATA_WIDTH)),
    5492 => std_logic_vector(to_unsigned(5420, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5493 => std_logic_vector(to_unsigned(6110, LDPC_TABLE_DATA_WIDTH)),
    5494 => std_logic_vector(to_unsigned(8551, LDPC_TABLE_DATA_WIDTH)),
    5495 => std_logic_vector(to_unsigned(1515, LDPC_TABLE_DATA_WIDTH)),
    5496 => std_logic_vector(to_unsigned(7404, LDPC_TABLE_DATA_WIDTH)),
    5497 => std_logic_vector(to_unsigned(4879, LDPC_TABLE_DATA_WIDTH)),
    5498 => std_logic_vector(to_unsigned(4946, LDPC_TABLE_DATA_WIDTH)),
    5499 => std_logic_vector(to_unsigned(5383, LDPC_TABLE_DATA_WIDTH)),
    5500 => std_logic_vector(to_unsigned(1831, LDPC_TABLE_DATA_WIDTH)),
    5501 => std_logic_vector(to_unsigned(3441, LDPC_TABLE_DATA_WIDTH)),
    5502 => std_logic_vector(to_unsigned(9569, LDPC_TABLE_DATA_WIDTH)),
    5503 => std_logic_vector(to_unsigned(10472, LDPC_TABLE_DATA_WIDTH)),
    5504 => std_logic_vector(to_unsigned(4306, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5505 => std_logic_vector(to_unsigned(1505, LDPC_TABLE_DATA_WIDTH)),
    5506 => std_logic_vector(to_unsigned(5682, LDPC_TABLE_DATA_WIDTH)),
    5507 => std_logic_vector(to_unsigned(7778, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5508 => std_logic_vector(to_unsigned(7172, LDPC_TABLE_DATA_WIDTH)),
    5509 => std_logic_vector(to_unsigned(6830, LDPC_TABLE_DATA_WIDTH)),
    5510 => std_logic_vector(to_unsigned(6623, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5511 => std_logic_vector(to_unsigned(7281, LDPC_TABLE_DATA_WIDTH)),
    5512 => std_logic_vector(to_unsigned(3941, LDPC_TABLE_DATA_WIDTH)),
    5513 => std_logic_vector(to_unsigned(3505, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5514 => std_logic_vector(to_unsigned(10270, LDPC_TABLE_DATA_WIDTH)),
    5515 => std_logic_vector(to_unsigned(8669, LDPC_TABLE_DATA_WIDTH)),
    5516 => std_logic_vector(to_unsigned(914, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5517 => std_logic_vector(to_unsigned(3622, LDPC_TABLE_DATA_WIDTH)),
    5518 => std_logic_vector(to_unsigned(7563, LDPC_TABLE_DATA_WIDTH)),
    5519 => std_logic_vector(to_unsigned(9388, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5520 => std_logic_vector(to_unsigned(9930, LDPC_TABLE_DATA_WIDTH)),
    5521 => std_logic_vector(to_unsigned(5058, LDPC_TABLE_DATA_WIDTH)),
    5522 => std_logic_vector(to_unsigned(4554, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5523 => std_logic_vector(to_unsigned(4844, LDPC_TABLE_DATA_WIDTH)),
    5524 => std_logic_vector(to_unsigned(9609, LDPC_TABLE_DATA_WIDTH)),
    5525 => std_logic_vector(to_unsigned(2707, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5526 => std_logic_vector(to_unsigned(6883, LDPC_TABLE_DATA_WIDTH)),
    5527 => std_logic_vector(to_unsigned(3237, LDPC_TABLE_DATA_WIDTH)),
    5528 => std_logic_vector(to_unsigned(1714, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5529 => std_logic_vector(to_unsigned(4768, LDPC_TABLE_DATA_WIDTH)),
    5530 => std_logic_vector(to_unsigned(3878, LDPC_TABLE_DATA_WIDTH)),
    5531 => std_logic_vector(to_unsigned(10017, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5532 => std_logic_vector(to_unsigned(10127, LDPC_TABLE_DATA_WIDTH)),
    5533 => std_logic_vector(to_unsigned(3334, LDPC_TABLE_DATA_WIDTH)),
    5534 => std_logic_vector(to_unsigned(8267, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C1_4
    5535 => std_logic_vector(to_unsigned(6295, LDPC_TABLE_DATA_WIDTH)),
    5536 => std_logic_vector(to_unsigned(9626, LDPC_TABLE_DATA_WIDTH)),
    5537 => std_logic_vector(to_unsigned(304, LDPC_TABLE_DATA_WIDTH)),
    5538 => std_logic_vector(to_unsigned(7695, LDPC_TABLE_DATA_WIDTH)),
    5539 => std_logic_vector(to_unsigned(4839, LDPC_TABLE_DATA_WIDTH)),
    5540 => std_logic_vector(to_unsigned(4936, LDPC_TABLE_DATA_WIDTH)),
    5541 => std_logic_vector(to_unsigned(1660, LDPC_TABLE_DATA_WIDTH)),
    5542 => std_logic_vector(to_unsigned(144, LDPC_TABLE_DATA_WIDTH)),
    5543 => std_logic_vector(to_unsigned(11203, LDPC_TABLE_DATA_WIDTH)),
    5544 => std_logic_vector(to_unsigned(5567, LDPC_TABLE_DATA_WIDTH)),
    5545 => std_logic_vector(to_unsigned(6347, LDPC_TABLE_DATA_WIDTH)),
    5546 => std_logic_vector(to_unsigned(12557, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5547 => std_logic_vector(to_unsigned(10691, LDPC_TABLE_DATA_WIDTH)),
    5548 => std_logic_vector(to_unsigned(4988, LDPC_TABLE_DATA_WIDTH)),
    5549 => std_logic_vector(to_unsigned(3859, LDPC_TABLE_DATA_WIDTH)),
    5550 => std_logic_vector(to_unsigned(3734, LDPC_TABLE_DATA_WIDTH)),
    5551 => std_logic_vector(to_unsigned(3071, LDPC_TABLE_DATA_WIDTH)),
    5552 => std_logic_vector(to_unsigned(3494, LDPC_TABLE_DATA_WIDTH)),
    5553 => std_logic_vector(to_unsigned(7687, LDPC_TABLE_DATA_WIDTH)),
    5554 => std_logic_vector(to_unsigned(10313, LDPC_TABLE_DATA_WIDTH)),
    5555 => std_logic_vector(to_unsigned(5964, LDPC_TABLE_DATA_WIDTH)),
    5556 => std_logic_vector(to_unsigned(8069, LDPC_TABLE_DATA_WIDTH)),
    5557 => std_logic_vector(to_unsigned(8296, LDPC_TABLE_DATA_WIDTH)),
    5558 => std_logic_vector(to_unsigned(11090, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5559 => std_logic_vector(to_unsigned(10774, LDPC_TABLE_DATA_WIDTH)),
    5560 => std_logic_vector(to_unsigned(3613, LDPC_TABLE_DATA_WIDTH)),
    5561 => std_logic_vector(to_unsigned(5208, LDPC_TABLE_DATA_WIDTH)),
    5562 => std_logic_vector(to_unsigned(11177, LDPC_TABLE_DATA_WIDTH)),
    5563 => std_logic_vector(to_unsigned(7676, LDPC_TABLE_DATA_WIDTH)),
    5564 => std_logic_vector(to_unsigned(3549, LDPC_TABLE_DATA_WIDTH)),
    5565 => std_logic_vector(to_unsigned(8746, LDPC_TABLE_DATA_WIDTH)),
    5566 => std_logic_vector(to_unsigned(6583, LDPC_TABLE_DATA_WIDTH)),
    5567 => std_logic_vector(to_unsigned(7239, LDPC_TABLE_DATA_WIDTH)),
    5568 => std_logic_vector(to_unsigned(12265, LDPC_TABLE_DATA_WIDTH)),
    5569 => std_logic_vector(to_unsigned(2674, LDPC_TABLE_DATA_WIDTH)),
    5570 => std_logic_vector(to_unsigned(4292, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5571 => std_logic_vector(to_unsigned(11869, LDPC_TABLE_DATA_WIDTH)),
    5572 => std_logic_vector(to_unsigned(3708, LDPC_TABLE_DATA_WIDTH)),
    5573 => std_logic_vector(to_unsigned(5981, LDPC_TABLE_DATA_WIDTH)),
    5574 => std_logic_vector(to_unsigned(8718, LDPC_TABLE_DATA_WIDTH)),
    5575 => std_logic_vector(to_unsigned(4908, LDPC_TABLE_DATA_WIDTH)),
    5576 => std_logic_vector(to_unsigned(10650, LDPC_TABLE_DATA_WIDTH)),
    5577 => std_logic_vector(to_unsigned(6805, LDPC_TABLE_DATA_WIDTH)),
    5578 => std_logic_vector(to_unsigned(3334, LDPC_TABLE_DATA_WIDTH)),
    5579 => std_logic_vector(to_unsigned(2627, LDPC_TABLE_DATA_WIDTH)),
    5580 => std_logic_vector(to_unsigned(10461, LDPC_TABLE_DATA_WIDTH)),
    5581 => std_logic_vector(to_unsigned(9285, LDPC_TABLE_DATA_WIDTH)),
    5582 => std_logic_vector(to_unsigned(11120, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5583 => std_logic_vector(to_unsigned(7844, LDPC_TABLE_DATA_WIDTH)),
    5584 => std_logic_vector(to_unsigned(3079, LDPC_TABLE_DATA_WIDTH)),
    5585 => std_logic_vector(to_unsigned(10773, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5586 => std_logic_vector(to_unsigned(3385, LDPC_TABLE_DATA_WIDTH)),
    5587 => std_logic_vector(to_unsigned(10854, LDPC_TABLE_DATA_WIDTH)),
    5588 => std_logic_vector(to_unsigned(5747, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5589 => std_logic_vector(to_unsigned(1360, LDPC_TABLE_DATA_WIDTH)),
    5590 => std_logic_vector(to_unsigned(12010, LDPC_TABLE_DATA_WIDTH)),
    5591 => std_logic_vector(to_unsigned(12202, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5592 => std_logic_vector(to_unsigned(6189, LDPC_TABLE_DATA_WIDTH)),
    5593 => std_logic_vector(to_unsigned(4241, LDPC_TABLE_DATA_WIDTH)),
    5594 => std_logic_vector(to_unsigned(2343, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5595 => std_logic_vector(to_unsigned(9840, LDPC_TABLE_DATA_WIDTH)),
    5596 => std_logic_vector(to_unsigned(12726, LDPC_TABLE_DATA_WIDTH)),
    5597 => std_logic_vector(to_unsigned(4977, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C2_3
    5598 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5599 => std_logic_vector(to_unsigned(2084, LDPC_TABLE_DATA_WIDTH)),
    5600 => std_logic_vector(to_unsigned(1613, LDPC_TABLE_DATA_WIDTH)),
    5601 => std_logic_vector(to_unsigned(1548, LDPC_TABLE_DATA_WIDTH)),
    5602 => std_logic_vector(to_unsigned(1286, LDPC_TABLE_DATA_WIDTH)),
    5603 => std_logic_vector(to_unsigned(1460, LDPC_TABLE_DATA_WIDTH)),
    5604 => std_logic_vector(to_unsigned(3196, LDPC_TABLE_DATA_WIDTH)),
    5605 => std_logic_vector(to_unsigned(4297, LDPC_TABLE_DATA_WIDTH)),
    5606 => std_logic_vector(to_unsigned(2481, LDPC_TABLE_DATA_WIDTH)),
    5607 => std_logic_vector(to_unsigned(3369, LDPC_TABLE_DATA_WIDTH)),
    5608 => std_logic_vector(to_unsigned(3451, LDPC_TABLE_DATA_WIDTH)),
    5609 => std_logic_vector(to_unsigned(4620, LDPC_TABLE_DATA_WIDTH)),
    5610 => std_logic_vector(to_unsigned(2622, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5611 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5612 => std_logic_vector(to_unsigned(122, LDPC_TABLE_DATA_WIDTH)),
    5613 => std_logic_vector(to_unsigned(1516, LDPC_TABLE_DATA_WIDTH)),
    5614 => std_logic_vector(to_unsigned(3448, LDPC_TABLE_DATA_WIDTH)),
    5615 => std_logic_vector(to_unsigned(2880, LDPC_TABLE_DATA_WIDTH)),
    5616 => std_logic_vector(to_unsigned(1407, LDPC_TABLE_DATA_WIDTH)),
    5617 => std_logic_vector(to_unsigned(1847, LDPC_TABLE_DATA_WIDTH)),
    5618 => std_logic_vector(to_unsigned(3799, LDPC_TABLE_DATA_WIDTH)),
    5619 => std_logic_vector(to_unsigned(3529, LDPC_TABLE_DATA_WIDTH)),
    5620 => std_logic_vector(to_unsigned(373, LDPC_TABLE_DATA_WIDTH)),
    5621 => std_logic_vector(to_unsigned(971, LDPC_TABLE_DATA_WIDTH)),
    5622 => std_logic_vector(to_unsigned(4358, LDPC_TABLE_DATA_WIDTH)),
    5623 => std_logic_vector(to_unsigned(3108, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5624 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5625 => std_logic_vector(to_unsigned(259, LDPC_TABLE_DATA_WIDTH)),
    5626 => std_logic_vector(to_unsigned(3399, LDPC_TABLE_DATA_WIDTH)),
    5627 => std_logic_vector(to_unsigned(929, LDPC_TABLE_DATA_WIDTH)),
    5628 => std_logic_vector(to_unsigned(2650, LDPC_TABLE_DATA_WIDTH)),
    5629 => std_logic_vector(to_unsigned(864, LDPC_TABLE_DATA_WIDTH)),
    5630 => std_logic_vector(to_unsigned(3996, LDPC_TABLE_DATA_WIDTH)),
    5631 => std_logic_vector(to_unsigned(3833, LDPC_TABLE_DATA_WIDTH)),
    5632 => std_logic_vector(to_unsigned(107, LDPC_TABLE_DATA_WIDTH)),
    5633 => std_logic_vector(to_unsigned(5287, LDPC_TABLE_DATA_WIDTH)),
    5634 => std_logic_vector(to_unsigned(164, LDPC_TABLE_DATA_WIDTH)),
    5635 => std_logic_vector(to_unsigned(3125, LDPC_TABLE_DATA_WIDTH)),
    5636 => std_logic_vector(to_unsigned(2350, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5637 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5638 => std_logic_vector(to_unsigned(342, LDPC_TABLE_DATA_WIDTH)),
    5639 => std_logic_vector(to_unsigned(3529, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5640 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5641 => std_logic_vector(to_unsigned(4198, LDPC_TABLE_DATA_WIDTH)),
    5642 => std_logic_vector(to_unsigned(2147, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5643 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5644 => std_logic_vector(to_unsigned(1880, LDPC_TABLE_DATA_WIDTH)),
    5645 => std_logic_vector(to_unsigned(4836, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5646 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5647 => std_logic_vector(to_unsigned(3864, LDPC_TABLE_DATA_WIDTH)),
    5648 => std_logic_vector(to_unsigned(4910, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5649 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5650 => std_logic_vector(to_unsigned(243, LDPC_TABLE_DATA_WIDTH)),
    5651 => std_logic_vector(to_unsigned(1542, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5652 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5653 => std_logic_vector(to_unsigned(3011, LDPC_TABLE_DATA_WIDTH)),
    5654 => std_logic_vector(to_unsigned(1436, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5655 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5656 => std_logic_vector(to_unsigned(2167, LDPC_TABLE_DATA_WIDTH)),
    5657 => std_logic_vector(to_unsigned(2512, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5658 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5659 => std_logic_vector(to_unsigned(4606, LDPC_TABLE_DATA_WIDTH)),
    5660 => std_logic_vector(to_unsigned(1003, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5661 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5662 => std_logic_vector(to_unsigned(2835, LDPC_TABLE_DATA_WIDTH)),
    5663 => std_logic_vector(to_unsigned(705, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5664 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5665 => std_logic_vector(to_unsigned(3426, LDPC_TABLE_DATA_WIDTH)),
    5666 => std_logic_vector(to_unsigned(2365, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5667 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5668 => std_logic_vector(to_unsigned(3848, LDPC_TABLE_DATA_WIDTH)),
    5669 => std_logic_vector(to_unsigned(2474, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5670 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5671 => std_logic_vector(to_unsigned(1360, LDPC_TABLE_DATA_WIDTH)),
    5672 => std_logic_vector(to_unsigned(1743, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5673 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5674 => std_logic_vector(to_unsigned(163, LDPC_TABLE_DATA_WIDTH)),
    5675 => std_logic_vector(to_unsigned(2536, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5676 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5677 => std_logic_vector(to_unsigned(2583, LDPC_TABLE_DATA_WIDTH)),
    5678 => std_logic_vector(to_unsigned(1180, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5679 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5680 => std_logic_vector(to_unsigned(1542, LDPC_TABLE_DATA_WIDTH)),
    5681 => std_logic_vector(to_unsigned(509, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5682 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5683 => std_logic_vector(to_unsigned(4418, LDPC_TABLE_DATA_WIDTH)),
    5684 => std_logic_vector(to_unsigned(1005, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5685 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5686 => std_logic_vector(to_unsigned(5212, LDPC_TABLE_DATA_WIDTH)),
    5687 => std_logic_vector(to_unsigned(5117, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5688 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5689 => std_logic_vector(to_unsigned(2155, LDPC_TABLE_DATA_WIDTH)),
    5690 => std_logic_vector(to_unsigned(2922, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5691 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5692 => std_logic_vector(to_unsigned(347, LDPC_TABLE_DATA_WIDTH)),
    5693 => std_logic_vector(to_unsigned(2696, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5694 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5695 => std_logic_vector(to_unsigned(226, LDPC_TABLE_DATA_WIDTH)),
    5696 => std_logic_vector(to_unsigned(4296, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5697 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5698 => std_logic_vector(to_unsigned(1560, LDPC_TABLE_DATA_WIDTH)),
    5699 => std_logic_vector(to_unsigned(487, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5700 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5701 => std_logic_vector(to_unsigned(3926, LDPC_TABLE_DATA_WIDTH)),
    5702 => std_logic_vector(to_unsigned(1640, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5703 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5704 => std_logic_vector(to_unsigned(149, LDPC_TABLE_DATA_WIDTH)),
    5705 => std_logic_vector(to_unsigned(2928, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5706 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5707 => std_logic_vector(to_unsigned(2364, LDPC_TABLE_DATA_WIDTH)),
    5708 => std_logic_vector(to_unsigned(563, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5709 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    5710 => std_logic_vector(to_unsigned(635, LDPC_TABLE_DATA_WIDTH)),
    5711 => std_logic_vector(to_unsigned(688, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5712 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    5713 => std_logic_vector(to_unsigned(231, LDPC_TABLE_DATA_WIDTH)),
    5714 => std_logic_vector(to_unsigned(1684, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5715 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    5716 => std_logic_vector(to_unsigned(1129, LDPC_TABLE_DATA_WIDTH)),
    5717 => std_logic_vector(to_unsigned(3894, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C2_5
    5718 => std_logic_vector(to_unsigned(5650, LDPC_TABLE_DATA_WIDTH)),
    5719 => std_logic_vector(to_unsigned(4143, LDPC_TABLE_DATA_WIDTH)),
    5720 => std_logic_vector(to_unsigned(8750, LDPC_TABLE_DATA_WIDTH)),
    5721 => std_logic_vector(to_unsigned(583, LDPC_TABLE_DATA_WIDTH)),
    5722 => std_logic_vector(to_unsigned(6720, LDPC_TABLE_DATA_WIDTH)),
    5723 => std_logic_vector(to_unsigned(8071, LDPC_TABLE_DATA_WIDTH)),
    5724 => std_logic_vector(to_unsigned(635, LDPC_TABLE_DATA_WIDTH)),
    5725 => std_logic_vector(to_unsigned(1767, LDPC_TABLE_DATA_WIDTH)),
    5726 => std_logic_vector(to_unsigned(1344, LDPC_TABLE_DATA_WIDTH)),
    5727 => std_logic_vector(to_unsigned(6922, LDPC_TABLE_DATA_WIDTH)),
    5728 => std_logic_vector(to_unsigned(738, LDPC_TABLE_DATA_WIDTH)),
    5729 => std_logic_vector(to_unsigned(6658, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5730 => std_logic_vector(to_unsigned(5696, LDPC_TABLE_DATA_WIDTH)),
    5731 => std_logic_vector(to_unsigned(1685, LDPC_TABLE_DATA_WIDTH)),
    5732 => std_logic_vector(to_unsigned(3207, LDPC_TABLE_DATA_WIDTH)),
    5733 => std_logic_vector(to_unsigned(415, LDPC_TABLE_DATA_WIDTH)),
    5734 => std_logic_vector(to_unsigned(7019, LDPC_TABLE_DATA_WIDTH)),
    5735 => std_logic_vector(to_unsigned(5023, LDPC_TABLE_DATA_WIDTH)),
    5736 => std_logic_vector(to_unsigned(5608, LDPC_TABLE_DATA_WIDTH)),
    5737 => std_logic_vector(to_unsigned(2605, LDPC_TABLE_DATA_WIDTH)),
    5738 => std_logic_vector(to_unsigned(857, LDPC_TABLE_DATA_WIDTH)),
    5739 => std_logic_vector(to_unsigned(6915, LDPC_TABLE_DATA_WIDTH)),
    5740 => std_logic_vector(to_unsigned(1770, LDPC_TABLE_DATA_WIDTH)),
    5741 => std_logic_vector(to_unsigned(8016, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5742 => std_logic_vector(to_unsigned(3992, LDPC_TABLE_DATA_WIDTH)),
    5743 => std_logic_vector(to_unsigned(771, LDPC_TABLE_DATA_WIDTH)),
    5744 => std_logic_vector(to_unsigned(2190, LDPC_TABLE_DATA_WIDTH)),
    5745 => std_logic_vector(to_unsigned(7258, LDPC_TABLE_DATA_WIDTH)),
    5746 => std_logic_vector(to_unsigned(8970, LDPC_TABLE_DATA_WIDTH)),
    5747 => std_logic_vector(to_unsigned(7792, LDPC_TABLE_DATA_WIDTH)),
    5748 => std_logic_vector(to_unsigned(1802, LDPC_TABLE_DATA_WIDTH)),
    5749 => std_logic_vector(to_unsigned(1866, LDPC_TABLE_DATA_WIDTH)),
    5750 => std_logic_vector(to_unsigned(6137, LDPC_TABLE_DATA_WIDTH)),
    5751 => std_logic_vector(to_unsigned(8841, LDPC_TABLE_DATA_WIDTH)),
    5752 => std_logic_vector(to_unsigned(886, LDPC_TABLE_DATA_WIDTH)),
    5753 => std_logic_vector(to_unsigned(1931, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5754 => std_logic_vector(to_unsigned(4108, LDPC_TABLE_DATA_WIDTH)),
    5755 => std_logic_vector(to_unsigned(3781, LDPC_TABLE_DATA_WIDTH)),
    5756 => std_logic_vector(to_unsigned(7577, LDPC_TABLE_DATA_WIDTH)),
    5757 => std_logic_vector(to_unsigned(6810, LDPC_TABLE_DATA_WIDTH)),
    5758 => std_logic_vector(to_unsigned(9322, LDPC_TABLE_DATA_WIDTH)),
    5759 => std_logic_vector(to_unsigned(8226, LDPC_TABLE_DATA_WIDTH)),
    5760 => std_logic_vector(to_unsigned(5396, LDPC_TABLE_DATA_WIDTH)),
    5761 => std_logic_vector(to_unsigned(5867, LDPC_TABLE_DATA_WIDTH)),
    5762 => std_logic_vector(to_unsigned(4428, LDPC_TABLE_DATA_WIDTH)),
    5763 => std_logic_vector(to_unsigned(8827, LDPC_TABLE_DATA_WIDTH)),
    5764 => std_logic_vector(to_unsigned(7766, LDPC_TABLE_DATA_WIDTH)),
    5765 => std_logic_vector(to_unsigned(2254, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5766 => std_logic_vector(to_unsigned(4247, LDPC_TABLE_DATA_WIDTH)),
    5767 => std_logic_vector(to_unsigned(888, LDPC_TABLE_DATA_WIDTH)),
    5768 => std_logic_vector(to_unsigned(4367, LDPC_TABLE_DATA_WIDTH)),
    5769 => std_logic_vector(to_unsigned(8821, LDPC_TABLE_DATA_WIDTH)),
    5770 => std_logic_vector(to_unsigned(9660, LDPC_TABLE_DATA_WIDTH)),
    5771 => std_logic_vector(to_unsigned(324, LDPC_TABLE_DATA_WIDTH)),
    5772 => std_logic_vector(to_unsigned(5864, LDPC_TABLE_DATA_WIDTH)),
    5773 => std_logic_vector(to_unsigned(4774, LDPC_TABLE_DATA_WIDTH)),
    5774 => std_logic_vector(to_unsigned(227, LDPC_TABLE_DATA_WIDTH)),
    5775 => std_logic_vector(to_unsigned(7889, LDPC_TABLE_DATA_WIDTH)),
    5776 => std_logic_vector(to_unsigned(6405, LDPC_TABLE_DATA_WIDTH)),
    5777 => std_logic_vector(to_unsigned(8963, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5778 => std_logic_vector(to_unsigned(9693, LDPC_TABLE_DATA_WIDTH)),
    5779 => std_logic_vector(to_unsigned(500, LDPC_TABLE_DATA_WIDTH)),
    5780 => std_logic_vector(to_unsigned(2520, LDPC_TABLE_DATA_WIDTH)),
    5781 => std_logic_vector(to_unsigned(2227, LDPC_TABLE_DATA_WIDTH)),
    5782 => std_logic_vector(to_unsigned(1811, LDPC_TABLE_DATA_WIDTH)),
    5783 => std_logic_vector(to_unsigned(9330, LDPC_TABLE_DATA_WIDTH)),
    5784 => std_logic_vector(to_unsigned(1928, LDPC_TABLE_DATA_WIDTH)),
    5785 => std_logic_vector(to_unsigned(5140, LDPC_TABLE_DATA_WIDTH)),
    5786 => std_logic_vector(to_unsigned(4030, LDPC_TABLE_DATA_WIDTH)),
    5787 => std_logic_vector(to_unsigned(4824, LDPC_TABLE_DATA_WIDTH)),
    5788 => std_logic_vector(to_unsigned(806, LDPC_TABLE_DATA_WIDTH)),
    5789 => std_logic_vector(to_unsigned(3134, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5790 => std_logic_vector(to_unsigned(1652, LDPC_TABLE_DATA_WIDTH)),
    5791 => std_logic_vector(to_unsigned(8171, LDPC_TABLE_DATA_WIDTH)),
    5792 => std_logic_vector(to_unsigned(1435, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5793 => std_logic_vector(to_unsigned(3366, LDPC_TABLE_DATA_WIDTH)),
    5794 => std_logic_vector(to_unsigned(6543, LDPC_TABLE_DATA_WIDTH)),
    5795 => std_logic_vector(to_unsigned(3745, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5796 => std_logic_vector(to_unsigned(9286, LDPC_TABLE_DATA_WIDTH)),
    5797 => std_logic_vector(to_unsigned(8509, LDPC_TABLE_DATA_WIDTH)),
    5798 => std_logic_vector(to_unsigned(4645, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5799 => std_logic_vector(to_unsigned(7397, LDPC_TABLE_DATA_WIDTH)),
    5800 => std_logic_vector(to_unsigned(5790, LDPC_TABLE_DATA_WIDTH)),
    5801 => std_logic_vector(to_unsigned(8972, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5802 => std_logic_vector(to_unsigned(6597, LDPC_TABLE_DATA_WIDTH)),
    5803 => std_logic_vector(to_unsigned(4422, LDPC_TABLE_DATA_WIDTH)),
    5804 => std_logic_vector(to_unsigned(1799, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5805 => std_logic_vector(to_unsigned(9276, LDPC_TABLE_DATA_WIDTH)),
    5806 => std_logic_vector(to_unsigned(4041, LDPC_TABLE_DATA_WIDTH)),
    5807 => std_logic_vector(to_unsigned(3847, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5808 => std_logic_vector(to_unsigned(8683, LDPC_TABLE_DATA_WIDTH)),
    5809 => std_logic_vector(to_unsigned(7378, LDPC_TABLE_DATA_WIDTH)),
    5810 => std_logic_vector(to_unsigned(4946, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5811 => std_logic_vector(to_unsigned(5348, LDPC_TABLE_DATA_WIDTH)),
    5812 => std_logic_vector(to_unsigned(1993, LDPC_TABLE_DATA_WIDTH)),
    5813 => std_logic_vector(to_unsigned(9186, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5814 => std_logic_vector(to_unsigned(6724, LDPC_TABLE_DATA_WIDTH)),
    5815 => std_logic_vector(to_unsigned(9015, LDPC_TABLE_DATA_WIDTH)),
    5816 => std_logic_vector(to_unsigned(5646, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5817 => std_logic_vector(to_unsigned(4502, LDPC_TABLE_DATA_WIDTH)),
    5818 => std_logic_vector(to_unsigned(4439, LDPC_TABLE_DATA_WIDTH)),
    5819 => std_logic_vector(to_unsigned(8474, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5820 => std_logic_vector(to_unsigned(5107, LDPC_TABLE_DATA_WIDTH)),
    5821 => std_logic_vector(to_unsigned(7342, LDPC_TABLE_DATA_WIDTH)),
    5822 => std_logic_vector(to_unsigned(9442, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5823 => std_logic_vector(to_unsigned(1387, LDPC_TABLE_DATA_WIDTH)),
    5824 => std_logic_vector(to_unsigned(8910, LDPC_TABLE_DATA_WIDTH)),
    5825 => std_logic_vector(to_unsigned(2660, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C3_4
    5826 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5827 => std_logic_vector(to_unsigned(3198, LDPC_TABLE_DATA_WIDTH)),
    5828 => std_logic_vector(to_unsigned(478, LDPC_TABLE_DATA_WIDTH)),
    5829 => std_logic_vector(to_unsigned(4207, LDPC_TABLE_DATA_WIDTH)),
    5830 => std_logic_vector(to_unsigned(1481, LDPC_TABLE_DATA_WIDTH)),
    5831 => std_logic_vector(to_unsigned(1009, LDPC_TABLE_DATA_WIDTH)),
    5832 => std_logic_vector(to_unsigned(2616, LDPC_TABLE_DATA_WIDTH)),
    5833 => std_logic_vector(to_unsigned(1924, LDPC_TABLE_DATA_WIDTH)),
    5834 => std_logic_vector(to_unsigned(3437, LDPC_TABLE_DATA_WIDTH)),
    5835 => std_logic_vector(to_unsigned(554, LDPC_TABLE_DATA_WIDTH)),
    5836 => std_logic_vector(to_unsigned(683, LDPC_TABLE_DATA_WIDTH)),
    5837 => std_logic_vector(to_unsigned(1801, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5838 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5839 => std_logic_vector(to_unsigned(2681, LDPC_TABLE_DATA_WIDTH)),
    5840 => std_logic_vector(to_unsigned(2135, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5841 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5842 => std_logic_vector(to_unsigned(3107, LDPC_TABLE_DATA_WIDTH)),
    5843 => std_logic_vector(to_unsigned(4027, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5844 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5845 => std_logic_vector(to_unsigned(2637, LDPC_TABLE_DATA_WIDTH)),
    5846 => std_logic_vector(to_unsigned(3373, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5847 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5848 => std_logic_vector(to_unsigned(3830, LDPC_TABLE_DATA_WIDTH)),
    5849 => std_logic_vector(to_unsigned(3449, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5850 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5851 => std_logic_vector(to_unsigned(4129, LDPC_TABLE_DATA_WIDTH)),
    5852 => std_logic_vector(to_unsigned(2060, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5853 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5854 => std_logic_vector(to_unsigned(4184, LDPC_TABLE_DATA_WIDTH)),
    5855 => std_logic_vector(to_unsigned(2742, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5856 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5857 => std_logic_vector(to_unsigned(3946, LDPC_TABLE_DATA_WIDTH)),
    5858 => std_logic_vector(to_unsigned(1070, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5859 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5860 => std_logic_vector(to_unsigned(2239, LDPC_TABLE_DATA_WIDTH)),
    5861 => std_logic_vector(to_unsigned(984, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5862 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5863 => std_logic_vector(to_unsigned(1458, LDPC_TABLE_DATA_WIDTH)),
    5864 => std_logic_vector(to_unsigned(3031, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5865 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5866 => std_logic_vector(to_unsigned(3003, LDPC_TABLE_DATA_WIDTH)),
    5867 => std_logic_vector(to_unsigned(1328, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5868 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5869 => std_logic_vector(to_unsigned(1137, LDPC_TABLE_DATA_WIDTH)),
    5870 => std_logic_vector(to_unsigned(1716, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5871 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5872 => std_logic_vector(to_unsigned(132, LDPC_TABLE_DATA_WIDTH)),
    5873 => std_logic_vector(to_unsigned(3725, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5874 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5875 => std_logic_vector(to_unsigned(1817, LDPC_TABLE_DATA_WIDTH)),
    5876 => std_logic_vector(to_unsigned(638, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5877 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5878 => std_logic_vector(to_unsigned(1774, LDPC_TABLE_DATA_WIDTH)),
    5879 => std_logic_vector(to_unsigned(3447, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5880 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5881 => std_logic_vector(to_unsigned(3632, LDPC_TABLE_DATA_WIDTH)),
    5882 => std_logic_vector(to_unsigned(1257, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5883 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5884 => std_logic_vector(to_unsigned(542, LDPC_TABLE_DATA_WIDTH)),
    5885 => std_logic_vector(to_unsigned(3694, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5886 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5887 => std_logic_vector(to_unsigned(1015, LDPC_TABLE_DATA_WIDTH)),
    5888 => std_logic_vector(to_unsigned(1945, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5889 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5890 => std_logic_vector(to_unsigned(1948, LDPC_TABLE_DATA_WIDTH)),
    5891 => std_logic_vector(to_unsigned(412, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5892 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5893 => std_logic_vector(to_unsigned(995, LDPC_TABLE_DATA_WIDTH)),
    5894 => std_logic_vector(to_unsigned(2238, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5895 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5896 => std_logic_vector(to_unsigned(4141, LDPC_TABLE_DATA_WIDTH)),
    5897 => std_logic_vector(to_unsigned(1907, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5898 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    5899 => std_logic_vector(to_unsigned(2480, LDPC_TABLE_DATA_WIDTH)),
    5900 => std_logic_vector(to_unsigned(3079, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5901 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    5902 => std_logic_vector(to_unsigned(3021, LDPC_TABLE_DATA_WIDTH)),
    5903 => std_logic_vector(to_unsigned(1088, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5904 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    5905 => std_logic_vector(to_unsigned(713, LDPC_TABLE_DATA_WIDTH)),
    5906 => std_logic_vector(to_unsigned(1379, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5907 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    5908 => std_logic_vector(to_unsigned(997, LDPC_TABLE_DATA_WIDTH)),
    5909 => std_logic_vector(to_unsigned(3903, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5910 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    5911 => std_logic_vector(to_unsigned(2323, LDPC_TABLE_DATA_WIDTH)),
    5912 => std_logic_vector(to_unsigned(3361, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5913 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    5914 => std_logic_vector(to_unsigned(1110, LDPC_TABLE_DATA_WIDTH)),
    5915 => std_logic_vector(to_unsigned(986, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5916 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    5917 => std_logic_vector(to_unsigned(2532, LDPC_TABLE_DATA_WIDTH)),
    5918 => std_logic_vector(to_unsigned(142, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5919 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    5920 => std_logic_vector(to_unsigned(1690, LDPC_TABLE_DATA_WIDTH)),
    5921 => std_logic_vector(to_unsigned(2405, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5922 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    5923 => std_logic_vector(to_unsigned(1298, LDPC_TABLE_DATA_WIDTH)),
    5924 => std_logic_vector(to_unsigned(1881, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5925 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    5926 => std_logic_vector(to_unsigned(615, LDPC_TABLE_DATA_WIDTH)),
    5927 => std_logic_vector(to_unsigned(174, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5928 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    5929 => std_logic_vector(to_unsigned(1648, LDPC_TABLE_DATA_WIDTH)),
    5930 => std_logic_vector(to_unsigned(3112, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5931 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    5932 => std_logic_vector(to_unsigned(1415, LDPC_TABLE_DATA_WIDTH)),
    5933 => std_logic_vector(to_unsigned(2808, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C3_5
    5934 => std_logic_vector(to_unsigned(2765, LDPC_TABLE_DATA_WIDTH)),
    5935 => std_logic_vector(to_unsigned(5713, LDPC_TABLE_DATA_WIDTH)),
    5936 => std_logic_vector(to_unsigned(6426, LDPC_TABLE_DATA_WIDTH)),
    5937 => std_logic_vector(to_unsigned(3596, LDPC_TABLE_DATA_WIDTH)),
    5938 => std_logic_vector(to_unsigned(1374, LDPC_TABLE_DATA_WIDTH)),
    5939 => std_logic_vector(to_unsigned(4811, LDPC_TABLE_DATA_WIDTH)),
    5940 => std_logic_vector(to_unsigned(2182, LDPC_TABLE_DATA_WIDTH)),
    5941 => std_logic_vector(to_unsigned(544, LDPC_TABLE_DATA_WIDTH)),
    5942 => std_logic_vector(to_unsigned(3394, LDPC_TABLE_DATA_WIDTH)),
    5943 => std_logic_vector(to_unsigned(2840, LDPC_TABLE_DATA_WIDTH)),
    5944 => std_logic_vector(to_unsigned(4310, LDPC_TABLE_DATA_WIDTH)),
    5945 => std_logic_vector(to_unsigned(771, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5946 => std_logic_vector(to_unsigned(4951, LDPC_TABLE_DATA_WIDTH)),
    5947 => std_logic_vector(to_unsigned(211, LDPC_TABLE_DATA_WIDTH)),
    5948 => std_logic_vector(to_unsigned(2208, LDPC_TABLE_DATA_WIDTH)),
    5949 => std_logic_vector(to_unsigned(723, LDPC_TABLE_DATA_WIDTH)),
    5950 => std_logic_vector(to_unsigned(1246, LDPC_TABLE_DATA_WIDTH)),
    5951 => std_logic_vector(to_unsigned(2928, LDPC_TABLE_DATA_WIDTH)),
    5952 => std_logic_vector(to_unsigned(398, LDPC_TABLE_DATA_WIDTH)),
    5953 => std_logic_vector(to_unsigned(5739, LDPC_TABLE_DATA_WIDTH)),
    5954 => std_logic_vector(to_unsigned(265, LDPC_TABLE_DATA_WIDTH)),
    5955 => std_logic_vector(to_unsigned(5601, LDPC_TABLE_DATA_WIDTH)),
    5956 => std_logic_vector(to_unsigned(5993, LDPC_TABLE_DATA_WIDTH)),
    5957 => std_logic_vector(to_unsigned(2615, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5958 => std_logic_vector(to_unsigned(210, LDPC_TABLE_DATA_WIDTH)),
    5959 => std_logic_vector(to_unsigned(4730, LDPC_TABLE_DATA_WIDTH)),
    5960 => std_logic_vector(to_unsigned(5777, LDPC_TABLE_DATA_WIDTH)),
    5961 => std_logic_vector(to_unsigned(3096, LDPC_TABLE_DATA_WIDTH)),
    5962 => std_logic_vector(to_unsigned(4282, LDPC_TABLE_DATA_WIDTH)),
    5963 => std_logic_vector(to_unsigned(6238, LDPC_TABLE_DATA_WIDTH)),
    5964 => std_logic_vector(to_unsigned(4939, LDPC_TABLE_DATA_WIDTH)),
    5965 => std_logic_vector(to_unsigned(1119, LDPC_TABLE_DATA_WIDTH)),
    5966 => std_logic_vector(to_unsigned(6463, LDPC_TABLE_DATA_WIDTH)),
    5967 => std_logic_vector(to_unsigned(5298, LDPC_TABLE_DATA_WIDTH)),
    5968 => std_logic_vector(to_unsigned(6320, LDPC_TABLE_DATA_WIDTH)),
    5969 => std_logic_vector(to_unsigned(4016, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5970 => std_logic_vector(to_unsigned(4167, LDPC_TABLE_DATA_WIDTH)),
    5971 => std_logic_vector(to_unsigned(2063, LDPC_TABLE_DATA_WIDTH)),
    5972 => std_logic_vector(to_unsigned(4757, LDPC_TABLE_DATA_WIDTH)),
    5973 => std_logic_vector(to_unsigned(3157, LDPC_TABLE_DATA_WIDTH)),
    5974 => std_logic_vector(to_unsigned(5664, LDPC_TABLE_DATA_WIDTH)),
    5975 => std_logic_vector(to_unsigned(3956, LDPC_TABLE_DATA_WIDTH)),
    5976 => std_logic_vector(to_unsigned(6045, LDPC_TABLE_DATA_WIDTH)),
    5977 => std_logic_vector(to_unsigned(563, LDPC_TABLE_DATA_WIDTH)),
    5978 => std_logic_vector(to_unsigned(4284, LDPC_TABLE_DATA_WIDTH)),
    5979 => std_logic_vector(to_unsigned(2441, LDPC_TABLE_DATA_WIDTH)),
    5980 => std_logic_vector(to_unsigned(3412, LDPC_TABLE_DATA_WIDTH)),
    5981 => std_logic_vector(to_unsigned(6334, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5982 => std_logic_vector(to_unsigned(4201, LDPC_TABLE_DATA_WIDTH)),
    5983 => std_logic_vector(to_unsigned(2428, LDPC_TABLE_DATA_WIDTH)),
    5984 => std_logic_vector(to_unsigned(4474, LDPC_TABLE_DATA_WIDTH)),
    5985 => std_logic_vector(to_unsigned(59, LDPC_TABLE_DATA_WIDTH)),
    5986 => std_logic_vector(to_unsigned(1721, LDPC_TABLE_DATA_WIDTH)),
    5987 => std_logic_vector(to_unsigned(736, LDPC_TABLE_DATA_WIDTH)),
    5988 => std_logic_vector(to_unsigned(2997, LDPC_TABLE_DATA_WIDTH)),
    5989 => std_logic_vector(to_unsigned(428, LDPC_TABLE_DATA_WIDTH)),
    5990 => std_logic_vector(to_unsigned(3807, LDPC_TABLE_DATA_WIDTH)),
    5991 => std_logic_vector(to_unsigned(1513, LDPC_TABLE_DATA_WIDTH)),
    5992 => std_logic_vector(to_unsigned(4732, LDPC_TABLE_DATA_WIDTH)),
    5993 => std_logic_vector(to_unsigned(6195, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    5994 => std_logic_vector(to_unsigned(2670, LDPC_TABLE_DATA_WIDTH)),
    5995 => std_logic_vector(to_unsigned(3081, LDPC_TABLE_DATA_WIDTH)),
    5996 => std_logic_vector(to_unsigned(5139, LDPC_TABLE_DATA_WIDTH)),
    5997 => std_logic_vector(to_unsigned(3736, LDPC_TABLE_DATA_WIDTH)),
    5998 => std_logic_vector(to_unsigned(1999, LDPC_TABLE_DATA_WIDTH)),
    5999 => std_logic_vector(to_unsigned(5889, LDPC_TABLE_DATA_WIDTH)),
    6000 => std_logic_vector(to_unsigned(4362, LDPC_TABLE_DATA_WIDTH)),
    6001 => std_logic_vector(to_unsigned(3806, LDPC_TABLE_DATA_WIDTH)),
    6002 => std_logic_vector(to_unsigned(4534, LDPC_TABLE_DATA_WIDTH)),
    6003 => std_logic_vector(to_unsigned(5409, LDPC_TABLE_DATA_WIDTH)),
    6004 => std_logic_vector(to_unsigned(6384, LDPC_TABLE_DATA_WIDTH)),
    6005 => std_logic_vector(to_unsigned(5809, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6006 => std_logic_vector(to_unsigned(5516, LDPC_TABLE_DATA_WIDTH)),
    6007 => std_logic_vector(to_unsigned(1622, LDPC_TABLE_DATA_WIDTH)),
    6008 => std_logic_vector(to_unsigned(2906, LDPC_TABLE_DATA_WIDTH)),
    6009 => std_logic_vector(to_unsigned(3285, LDPC_TABLE_DATA_WIDTH)),
    6010 => std_logic_vector(to_unsigned(1257, LDPC_TABLE_DATA_WIDTH)),
    6011 => std_logic_vector(to_unsigned(5797, LDPC_TABLE_DATA_WIDTH)),
    6012 => std_logic_vector(to_unsigned(3816, LDPC_TABLE_DATA_WIDTH)),
    6013 => std_logic_vector(to_unsigned(817, LDPC_TABLE_DATA_WIDTH)),
    6014 => std_logic_vector(to_unsigned(875, LDPC_TABLE_DATA_WIDTH)),
    6015 => std_logic_vector(to_unsigned(2311, LDPC_TABLE_DATA_WIDTH)),
    6016 => std_logic_vector(to_unsigned(3543, LDPC_TABLE_DATA_WIDTH)),
    6017 => std_logic_vector(to_unsigned(1205, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6018 => std_logic_vector(to_unsigned(4244, LDPC_TABLE_DATA_WIDTH)),
    6019 => std_logic_vector(to_unsigned(2184, LDPC_TABLE_DATA_WIDTH)),
    6020 => std_logic_vector(to_unsigned(5415, LDPC_TABLE_DATA_WIDTH)),
    6021 => std_logic_vector(to_unsigned(1705, LDPC_TABLE_DATA_WIDTH)),
    6022 => std_logic_vector(to_unsigned(5642, LDPC_TABLE_DATA_WIDTH)),
    6023 => std_logic_vector(to_unsigned(4886, LDPC_TABLE_DATA_WIDTH)),
    6024 => std_logic_vector(to_unsigned(2333, LDPC_TABLE_DATA_WIDTH)),
    6025 => std_logic_vector(to_unsigned(287, LDPC_TABLE_DATA_WIDTH)),
    6026 => std_logic_vector(to_unsigned(1848, LDPC_TABLE_DATA_WIDTH)),
    6027 => std_logic_vector(to_unsigned(1121, LDPC_TABLE_DATA_WIDTH)),
    6028 => std_logic_vector(to_unsigned(3595, LDPC_TABLE_DATA_WIDTH)),
    6029 => std_logic_vector(to_unsigned(6022, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6030 => std_logic_vector(to_unsigned(2142, LDPC_TABLE_DATA_WIDTH)),
    6031 => std_logic_vector(to_unsigned(2830, LDPC_TABLE_DATA_WIDTH)),
    6032 => std_logic_vector(to_unsigned(4069, LDPC_TABLE_DATA_WIDTH)),
    6033 => std_logic_vector(to_unsigned(5654, LDPC_TABLE_DATA_WIDTH)),
    6034 => std_logic_vector(to_unsigned(1295, LDPC_TABLE_DATA_WIDTH)),
    6035 => std_logic_vector(to_unsigned(2951, LDPC_TABLE_DATA_WIDTH)),
    6036 => std_logic_vector(to_unsigned(3919, LDPC_TABLE_DATA_WIDTH)),
    6037 => std_logic_vector(to_unsigned(1356, LDPC_TABLE_DATA_WIDTH)),
    6038 => std_logic_vector(to_unsigned(884, LDPC_TABLE_DATA_WIDTH)),
    6039 => std_logic_vector(to_unsigned(1786, LDPC_TABLE_DATA_WIDTH)),
    6040 => std_logic_vector(to_unsigned(396, LDPC_TABLE_DATA_WIDTH)),
    6041 => std_logic_vector(to_unsigned(4738, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6042 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6043 => std_logic_vector(to_unsigned(2161, LDPC_TABLE_DATA_WIDTH)),
    6044 => std_logic_vector(to_unsigned(2653, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6045 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6046 => std_logic_vector(to_unsigned(1380, LDPC_TABLE_DATA_WIDTH)),
    6047 => std_logic_vector(to_unsigned(1461, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6048 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6049 => std_logic_vector(to_unsigned(2502, LDPC_TABLE_DATA_WIDTH)),
    6050 => std_logic_vector(to_unsigned(3707, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6051 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6052 => std_logic_vector(to_unsigned(3971, LDPC_TABLE_DATA_WIDTH)),
    6053 => std_logic_vector(to_unsigned(1057, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6054 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6055 => std_logic_vector(to_unsigned(5985, LDPC_TABLE_DATA_WIDTH)),
    6056 => std_logic_vector(to_unsigned(6062, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6057 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6058 => std_logic_vector(to_unsigned(1733, LDPC_TABLE_DATA_WIDTH)),
    6059 => std_logic_vector(to_unsigned(6028, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6060 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6061 => std_logic_vector(to_unsigned(3786, LDPC_TABLE_DATA_WIDTH)),
    6062 => std_logic_vector(to_unsigned(1936, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6063 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6064 => std_logic_vector(to_unsigned(4292, LDPC_TABLE_DATA_WIDTH)),
    6065 => std_logic_vector(to_unsigned(956, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6066 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    6067 => std_logic_vector(to_unsigned(5692, LDPC_TABLE_DATA_WIDTH)),
    6068 => std_logic_vector(to_unsigned(3417, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6069 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    6070 => std_logic_vector(to_unsigned(266, LDPC_TABLE_DATA_WIDTH)),
    6071 => std_logic_vector(to_unsigned(4878, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6072 => std_logic_vector(to_unsigned(10, LDPC_TABLE_DATA_WIDTH)),
    6073 => std_logic_vector(to_unsigned(4913, LDPC_TABLE_DATA_WIDTH)),
    6074 => std_logic_vector(to_unsigned(3247, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6075 => std_logic_vector(to_unsigned(11, LDPC_TABLE_DATA_WIDTH)),
    6076 => std_logic_vector(to_unsigned(4763, LDPC_TABLE_DATA_WIDTH)),
    6077 => std_logic_vector(to_unsigned(3937, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6078 => std_logic_vector(to_unsigned(12, LDPC_TABLE_DATA_WIDTH)),
    6079 => std_logic_vector(to_unsigned(3590, LDPC_TABLE_DATA_WIDTH)),
    6080 => std_logic_vector(to_unsigned(2903, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6081 => std_logic_vector(to_unsigned(13, LDPC_TABLE_DATA_WIDTH)),
    6082 => std_logic_vector(to_unsigned(2566, LDPC_TABLE_DATA_WIDTH)),
    6083 => std_logic_vector(to_unsigned(4215, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6084 => std_logic_vector(to_unsigned(14, LDPC_TABLE_DATA_WIDTH)),
    6085 => std_logic_vector(to_unsigned(5208, LDPC_TABLE_DATA_WIDTH)),
    6086 => std_logic_vector(to_unsigned(4707, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6087 => std_logic_vector(to_unsigned(15, LDPC_TABLE_DATA_WIDTH)),
    6088 => std_logic_vector(to_unsigned(3940, LDPC_TABLE_DATA_WIDTH)),
    6089 => std_logic_vector(to_unsigned(3388, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6090 => std_logic_vector(to_unsigned(16, LDPC_TABLE_DATA_WIDTH)),
    6091 => std_logic_vector(to_unsigned(5109, LDPC_TABLE_DATA_WIDTH)),
    6092 => std_logic_vector(to_unsigned(4556, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6093 => std_logic_vector(to_unsigned(17, LDPC_TABLE_DATA_WIDTH)),
    6094 => std_logic_vector(to_unsigned(4908, LDPC_TABLE_DATA_WIDTH)),
    6095 => std_logic_vector(to_unsigned(4177, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C4_5
    6096 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6097 => std_logic_vector(to_unsigned(896, LDPC_TABLE_DATA_WIDTH)),
    6098 => std_logic_vector(to_unsigned(1565, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6099 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6100 => std_logic_vector(to_unsigned(2493, LDPC_TABLE_DATA_WIDTH)),
    6101 => std_logic_vector(to_unsigned(184, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6102 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6103 => std_logic_vector(to_unsigned(212, LDPC_TABLE_DATA_WIDTH)),
    6104 => std_logic_vector(to_unsigned(3210, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6105 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    6106 => std_logic_vector(to_unsigned(727, LDPC_TABLE_DATA_WIDTH)),
    6107 => std_logic_vector(to_unsigned(1339, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6108 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    6109 => std_logic_vector(to_unsigned(3428, LDPC_TABLE_DATA_WIDTH)),
    6110 => std_logic_vector(to_unsigned(612, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6111 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6112 => std_logic_vector(to_unsigned(2663, LDPC_TABLE_DATA_WIDTH)),
    6113 => std_logic_vector(to_unsigned(1947, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6114 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6115 => std_logic_vector(to_unsigned(230, LDPC_TABLE_DATA_WIDTH)),
    6116 => std_logic_vector(to_unsigned(2695, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6117 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6118 => std_logic_vector(to_unsigned(2025, LDPC_TABLE_DATA_WIDTH)),
    6119 => std_logic_vector(to_unsigned(2794, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6120 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6121 => std_logic_vector(to_unsigned(3039, LDPC_TABLE_DATA_WIDTH)),
    6122 => std_logic_vector(to_unsigned(283, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6123 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6124 => std_logic_vector(to_unsigned(862, LDPC_TABLE_DATA_WIDTH)),
    6125 => std_logic_vector(to_unsigned(2889, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6126 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6127 => std_logic_vector(to_unsigned(376, LDPC_TABLE_DATA_WIDTH)),
    6128 => std_logic_vector(to_unsigned(2110, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6129 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6130 => std_logic_vector(to_unsigned(2034, LDPC_TABLE_DATA_WIDTH)),
    6131 => std_logic_vector(to_unsigned(2286, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6132 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6133 => std_logic_vector(to_unsigned(951, LDPC_TABLE_DATA_WIDTH)),
    6134 => std_logic_vector(to_unsigned(2068, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6135 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    6136 => std_logic_vector(to_unsigned(3108, LDPC_TABLE_DATA_WIDTH)),
    6137 => std_logic_vector(to_unsigned(3542, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6138 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    6139 => std_logic_vector(to_unsigned(307, LDPC_TABLE_DATA_WIDTH)),
    6140 => std_logic_vector(to_unsigned(1421, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6141 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6142 => std_logic_vector(to_unsigned(2272, LDPC_TABLE_DATA_WIDTH)),
    6143 => std_logic_vector(to_unsigned(1197, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6144 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6145 => std_logic_vector(to_unsigned(1800, LDPC_TABLE_DATA_WIDTH)),
    6146 => std_logic_vector(to_unsigned(3280, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6147 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6148 => std_logic_vector(to_unsigned(331, LDPC_TABLE_DATA_WIDTH)),
    6149 => std_logic_vector(to_unsigned(2308, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6150 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6151 => std_logic_vector(to_unsigned(465, LDPC_TABLE_DATA_WIDTH)),
    6152 => std_logic_vector(to_unsigned(2552, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6153 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6154 => std_logic_vector(to_unsigned(1038, LDPC_TABLE_DATA_WIDTH)),
    6155 => std_logic_vector(to_unsigned(2479, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6156 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6157 => std_logic_vector(to_unsigned(1383, LDPC_TABLE_DATA_WIDTH)),
    6158 => std_logic_vector(to_unsigned(343, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6159 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6160 => std_logic_vector(to_unsigned(94, LDPC_TABLE_DATA_WIDTH)),
    6161 => std_logic_vector(to_unsigned(236, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6162 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6163 => std_logic_vector(to_unsigned(2619, LDPC_TABLE_DATA_WIDTH)),
    6164 => std_logic_vector(to_unsigned(121, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6165 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    6166 => std_logic_vector(to_unsigned(1497, LDPC_TABLE_DATA_WIDTH)),
    6167 => std_logic_vector(to_unsigned(2774, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6168 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    6169 => std_logic_vector(to_unsigned(2116, LDPC_TABLE_DATA_WIDTH)),
    6170 => std_logic_vector(to_unsigned(1855, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6171 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6172 => std_logic_vector(to_unsigned(722, LDPC_TABLE_DATA_WIDTH)),
    6173 => std_logic_vector(to_unsigned(1584, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6174 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6175 => std_logic_vector(to_unsigned(2767, LDPC_TABLE_DATA_WIDTH)),
    6176 => std_logic_vector(to_unsigned(1881, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6177 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6178 => std_logic_vector(to_unsigned(2701, LDPC_TABLE_DATA_WIDTH)),
    6179 => std_logic_vector(to_unsigned(1610, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6180 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6181 => std_logic_vector(to_unsigned(3283, LDPC_TABLE_DATA_WIDTH)),
    6182 => std_logic_vector(to_unsigned(1732, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6183 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6184 => std_logic_vector(to_unsigned(168, LDPC_TABLE_DATA_WIDTH)),
    6185 => std_logic_vector(to_unsigned(1099, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6186 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6187 => std_logic_vector(to_unsigned(3074, LDPC_TABLE_DATA_WIDTH)),
    6188 => std_logic_vector(to_unsigned(243, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6189 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6190 => std_logic_vector(to_unsigned(3460, LDPC_TABLE_DATA_WIDTH)),
    6191 => std_logic_vector(to_unsigned(945, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6192 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6193 => std_logic_vector(to_unsigned(2049, LDPC_TABLE_DATA_WIDTH)),
    6194 => std_logic_vector(to_unsigned(1746, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6195 => std_logic_vector(to_unsigned(8, LDPC_TABLE_DATA_WIDTH)),
    6196 => std_logic_vector(to_unsigned(566, LDPC_TABLE_DATA_WIDTH)),
    6197 => std_logic_vector(to_unsigned(1427, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6198 => std_logic_vector(to_unsigned(9, LDPC_TABLE_DATA_WIDTH)),
    6199 => std_logic_vector(to_unsigned(3545, LDPC_TABLE_DATA_WIDTH)),
    6200 => std_logic_vector(to_unsigned(1168, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C5_6
    6201 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6202 => std_logic_vector(to_unsigned(2409, LDPC_TABLE_DATA_WIDTH)),
    6203 => std_logic_vector(to_unsigned(499, LDPC_TABLE_DATA_WIDTH)),
    6204 => std_logic_vector(to_unsigned(1481, LDPC_TABLE_DATA_WIDTH)),
    6205 => std_logic_vector(to_unsigned(908, LDPC_TABLE_DATA_WIDTH)),
    6206 => std_logic_vector(to_unsigned(559, LDPC_TABLE_DATA_WIDTH)),
    6207 => std_logic_vector(to_unsigned(716, LDPC_TABLE_DATA_WIDTH)),
    6208 => std_logic_vector(to_unsigned(1270, LDPC_TABLE_DATA_WIDTH)),
    6209 => std_logic_vector(to_unsigned(333, LDPC_TABLE_DATA_WIDTH)),
    6210 => std_logic_vector(to_unsigned(2508, LDPC_TABLE_DATA_WIDTH)),
    6211 => std_logic_vector(to_unsigned(2264, LDPC_TABLE_DATA_WIDTH)),
    6212 => std_logic_vector(to_unsigned(1702, LDPC_TABLE_DATA_WIDTH)),
    6213 => std_logic_vector(to_unsigned(2805, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6214 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6215 => std_logic_vector(to_unsigned(2447, LDPC_TABLE_DATA_WIDTH)),
    6216 => std_logic_vector(to_unsigned(1926, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6217 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6218 => std_logic_vector(to_unsigned(414, LDPC_TABLE_DATA_WIDTH)),
    6219 => std_logic_vector(to_unsigned(1224, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6220 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6221 => std_logic_vector(to_unsigned(2114, LDPC_TABLE_DATA_WIDTH)),
    6222 => std_logic_vector(to_unsigned(842, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6223 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6224 => std_logic_vector(to_unsigned(212, LDPC_TABLE_DATA_WIDTH)),
    6225 => std_logic_vector(to_unsigned(573, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6226 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6227 => std_logic_vector(to_unsigned(2383, LDPC_TABLE_DATA_WIDTH)),
    6228 => std_logic_vector(to_unsigned(2112, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6229 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6230 => std_logic_vector(to_unsigned(2286, LDPC_TABLE_DATA_WIDTH)),
    6231 => std_logic_vector(to_unsigned(2348, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6232 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6233 => std_logic_vector(to_unsigned(545, LDPC_TABLE_DATA_WIDTH)),
    6234 => std_logic_vector(to_unsigned(819, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6235 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6236 => std_logic_vector(to_unsigned(1264, LDPC_TABLE_DATA_WIDTH)),
    6237 => std_logic_vector(to_unsigned(143, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6238 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6239 => std_logic_vector(to_unsigned(1701, LDPC_TABLE_DATA_WIDTH)),
    6240 => std_logic_vector(to_unsigned(2258, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6241 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6242 => std_logic_vector(to_unsigned(964, LDPC_TABLE_DATA_WIDTH)),
    6243 => std_logic_vector(to_unsigned(166, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6244 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6245 => std_logic_vector(to_unsigned(114, LDPC_TABLE_DATA_WIDTH)),
    6246 => std_logic_vector(to_unsigned(2413, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6247 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6248 => std_logic_vector(to_unsigned(2243, LDPC_TABLE_DATA_WIDTH)),
    6249 => std_logic_vector(to_unsigned(81, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6250 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6251 => std_logic_vector(to_unsigned(1245, LDPC_TABLE_DATA_WIDTH)),
    6252 => std_logic_vector(to_unsigned(1581, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6253 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6254 => std_logic_vector(to_unsigned(775, LDPC_TABLE_DATA_WIDTH)),
    6255 => std_logic_vector(to_unsigned(169, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6256 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6257 => std_logic_vector(to_unsigned(1696, LDPC_TABLE_DATA_WIDTH)),
    6258 => std_logic_vector(to_unsigned(1104, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6259 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6260 => std_logic_vector(to_unsigned(1914, LDPC_TABLE_DATA_WIDTH)),
    6261 => std_logic_vector(to_unsigned(2831, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6262 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6263 => std_logic_vector(to_unsigned(532, LDPC_TABLE_DATA_WIDTH)),
    6264 => std_logic_vector(to_unsigned(1450, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6265 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6266 => std_logic_vector(to_unsigned(91, LDPC_TABLE_DATA_WIDTH)),
    6267 => std_logic_vector(to_unsigned(974, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6268 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6269 => std_logic_vector(to_unsigned(497, LDPC_TABLE_DATA_WIDTH)),
    6270 => std_logic_vector(to_unsigned(2228, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6271 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6272 => std_logic_vector(to_unsigned(2326, LDPC_TABLE_DATA_WIDTH)),
    6273 => std_logic_vector(to_unsigned(1579, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6274 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6275 => std_logic_vector(to_unsigned(2482, LDPC_TABLE_DATA_WIDTH)),
    6276 => std_logic_vector(to_unsigned(256, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6277 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6278 => std_logic_vector(to_unsigned(1117, LDPC_TABLE_DATA_WIDTH)),
    6279 => std_logic_vector(to_unsigned(1261, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6280 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6281 => std_logic_vector(to_unsigned(1257, LDPC_TABLE_DATA_WIDTH)),
    6282 => std_logic_vector(to_unsigned(1658, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6283 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6284 => std_logic_vector(to_unsigned(1478, LDPC_TABLE_DATA_WIDTH)),
    6285 => std_logic_vector(to_unsigned(1225, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6286 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6287 => std_logic_vector(to_unsigned(2511, LDPC_TABLE_DATA_WIDTH)),
    6288 => std_logic_vector(to_unsigned(980, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6289 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6290 => std_logic_vector(to_unsigned(2320, LDPC_TABLE_DATA_WIDTH)),
    6291 => std_logic_vector(to_unsigned(2675, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6292 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6293 => std_logic_vector(to_unsigned(435, LDPC_TABLE_DATA_WIDTH)),
    6294 => std_logic_vector(to_unsigned(1278, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6295 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6296 => std_logic_vector(to_unsigned(228, LDPC_TABLE_DATA_WIDTH)),
    6297 => std_logic_vector(to_unsigned(503, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6298 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6299 => std_logic_vector(to_unsigned(1885, LDPC_TABLE_DATA_WIDTH)),
    6300 => std_logic_vector(to_unsigned(2369, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6301 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6302 => std_logic_vector(to_unsigned(57, LDPC_TABLE_DATA_WIDTH)),
    6303 => std_logic_vector(to_unsigned(483, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6304 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6305 => std_logic_vector(to_unsigned(838, LDPC_TABLE_DATA_WIDTH)),
    6306 => std_logic_vector(to_unsigned(1050, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6307 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6308 => std_logic_vector(to_unsigned(1231, LDPC_TABLE_DATA_WIDTH)),
    6309 => std_logic_vector(to_unsigned(1990, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6310 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6311 => std_logic_vector(to_unsigned(1738, LDPC_TABLE_DATA_WIDTH)),
    6312 => std_logic_vector(to_unsigned(68, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6313 => std_logic_vector(to_unsigned(5, LDPC_TABLE_DATA_WIDTH)),
    6314 => std_logic_vector(to_unsigned(2392, LDPC_TABLE_DATA_WIDTH)),
    6315 => std_logic_vector(to_unsigned(951, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6316 => std_logic_vector(to_unsigned(6, LDPC_TABLE_DATA_WIDTH)),
    6317 => std_logic_vector(to_unsigned(163, LDPC_TABLE_DATA_WIDTH)),
    6318 => std_logic_vector(to_unsigned(645, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6319 => std_logic_vector(to_unsigned(7, LDPC_TABLE_DATA_WIDTH)),
    6320 => std_logic_vector(to_unsigned(2644, LDPC_TABLE_DATA_WIDTH)),
    6321 => std_logic_vector(to_unsigned(1704, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    -- Table for fecframe_short, C8_9
    6322 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6323 => std_logic_vector(to_unsigned(1558, LDPC_TABLE_DATA_WIDTH)),
    6324 => std_logic_vector(to_unsigned(712, LDPC_TABLE_DATA_WIDTH)),
    6325 => std_logic_vector(to_unsigned(805, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6326 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6327 => std_logic_vector(to_unsigned(1450, LDPC_TABLE_DATA_WIDTH)),
    6328 => std_logic_vector(to_unsigned(873, LDPC_TABLE_DATA_WIDTH)),
    6329 => std_logic_vector(to_unsigned(1337, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6330 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6331 => std_logic_vector(to_unsigned(1741, LDPC_TABLE_DATA_WIDTH)),
    6332 => std_logic_vector(to_unsigned(1129, LDPC_TABLE_DATA_WIDTH)),
    6333 => std_logic_vector(to_unsigned(1184, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6334 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6335 => std_logic_vector(to_unsigned(294, LDPC_TABLE_DATA_WIDTH)),
    6336 => std_logic_vector(to_unsigned(806, LDPC_TABLE_DATA_WIDTH)),
    6337 => std_logic_vector(to_unsigned(1566, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6338 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6339 => std_logic_vector(to_unsigned(482, LDPC_TABLE_DATA_WIDTH)),
    6340 => std_logic_vector(to_unsigned(605, LDPC_TABLE_DATA_WIDTH)),
    6341 => std_logic_vector(to_unsigned(923, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6342 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6343 => std_logic_vector(to_unsigned(926, LDPC_TABLE_DATA_WIDTH)),
    6344 => std_logic_vector(to_unsigned(1578, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6345 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6346 => std_logic_vector(to_unsigned(777, LDPC_TABLE_DATA_WIDTH)),
    6347 => std_logic_vector(to_unsigned(1374, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6348 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6349 => std_logic_vector(to_unsigned(608, LDPC_TABLE_DATA_WIDTH)),
    6350 => std_logic_vector(to_unsigned(151, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6351 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6352 => std_logic_vector(to_unsigned(1195, LDPC_TABLE_DATA_WIDTH)),
    6353 => std_logic_vector(to_unsigned(210, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6354 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6355 => std_logic_vector(to_unsigned(1484, LDPC_TABLE_DATA_WIDTH)),
    6356 => std_logic_vector(to_unsigned(692, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6357 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6358 => std_logic_vector(to_unsigned(427, LDPC_TABLE_DATA_WIDTH)),
    6359 => std_logic_vector(to_unsigned(488, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6360 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6361 => std_logic_vector(to_unsigned(828, LDPC_TABLE_DATA_WIDTH)),
    6362 => std_logic_vector(to_unsigned(1124, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6363 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6364 => std_logic_vector(to_unsigned(874, LDPC_TABLE_DATA_WIDTH)),
    6365 => std_logic_vector(to_unsigned(1366, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6366 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6367 => std_logic_vector(to_unsigned(1500, LDPC_TABLE_DATA_WIDTH)),
    6368 => std_logic_vector(to_unsigned(835, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6369 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6370 => std_logic_vector(to_unsigned(1496, LDPC_TABLE_DATA_WIDTH)),
    6371 => std_logic_vector(to_unsigned(502, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6372 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6373 => std_logic_vector(to_unsigned(1006, LDPC_TABLE_DATA_WIDTH)),
    6374 => std_logic_vector(to_unsigned(1701, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6375 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6376 => std_logic_vector(to_unsigned(1155, LDPC_TABLE_DATA_WIDTH)),
    6377 => std_logic_vector(to_unsigned(97, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6378 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6379 => std_logic_vector(to_unsigned(657, LDPC_TABLE_DATA_WIDTH)),
    6380 => std_logic_vector(to_unsigned(1403, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6381 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6382 => std_logic_vector(to_unsigned(1453, LDPC_TABLE_DATA_WIDTH)),
    6383 => std_logic_vector(to_unsigned(624, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6384 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6385 => std_logic_vector(to_unsigned(429, LDPC_TABLE_DATA_WIDTH)),
    6386 => std_logic_vector(to_unsigned(1495, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6387 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6388 => std_logic_vector(to_unsigned(809, LDPC_TABLE_DATA_WIDTH)),
    6389 => std_logic_vector(to_unsigned(385, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6390 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6391 => std_logic_vector(to_unsigned(367, LDPC_TABLE_DATA_WIDTH)),
    6392 => std_logic_vector(to_unsigned(151, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6393 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6394 => std_logic_vector(to_unsigned(1323, LDPC_TABLE_DATA_WIDTH)),
    6395 => std_logic_vector(to_unsigned(202, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6396 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6397 => std_logic_vector(to_unsigned(960, LDPC_TABLE_DATA_WIDTH)),
    6398 => std_logic_vector(to_unsigned(318, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6399 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6400 => std_logic_vector(to_unsigned(1451, LDPC_TABLE_DATA_WIDTH)),
    6401 => std_logic_vector(to_unsigned(1039, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6402 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6403 => std_logic_vector(to_unsigned(1098, LDPC_TABLE_DATA_WIDTH)),
    6404 => std_logic_vector(to_unsigned(1722, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6405 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6406 => std_logic_vector(to_unsigned(1015, LDPC_TABLE_DATA_WIDTH)),
    6407 => std_logic_vector(to_unsigned(1428, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6408 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6409 => std_logic_vector(to_unsigned(1261, LDPC_TABLE_DATA_WIDTH)),
    6410 => std_logic_vector(to_unsigned(1564, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6411 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6412 => std_logic_vector(to_unsigned(544, LDPC_TABLE_DATA_WIDTH)),
    6413 => std_logic_vector(to_unsigned(1190, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6414 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6415 => std_logic_vector(to_unsigned(1472, LDPC_TABLE_DATA_WIDTH)),
    6416 => std_logic_vector(to_unsigned(1246, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6417 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6418 => std_logic_vector(to_unsigned(508, LDPC_TABLE_DATA_WIDTH)),
    6419 => std_logic_vector(to_unsigned(630, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6420 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6421 => std_logic_vector(to_unsigned(421, LDPC_TABLE_DATA_WIDTH)),
    6422 => std_logic_vector(to_unsigned(1704, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6423 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6424 => std_logic_vector(to_unsigned(284, LDPC_TABLE_DATA_WIDTH)),
    6425 => std_logic_vector(to_unsigned(898, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6426 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6427 => std_logic_vector(to_unsigned(392, LDPC_TABLE_DATA_WIDTH)),
    6428 => std_logic_vector(to_unsigned(577, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6429 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6430 => std_logic_vector(to_unsigned(1155, LDPC_TABLE_DATA_WIDTH)),
    6431 => std_logic_vector(to_unsigned(556, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6432 => std_logic_vector(to_unsigned(0, LDPC_TABLE_DATA_WIDTH)),
    6433 => std_logic_vector(to_unsigned(631, LDPC_TABLE_DATA_WIDTH)),
    6434 => std_logic_vector(to_unsigned(1000, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6435 => std_logic_vector(to_unsigned(1, LDPC_TABLE_DATA_WIDTH)),
    6436 => std_logic_vector(to_unsigned(732, LDPC_TABLE_DATA_WIDTH)),
    6437 => std_logic_vector(to_unsigned(1368, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6438 => std_logic_vector(to_unsigned(2, LDPC_TABLE_DATA_WIDTH)),
    6439 => std_logic_vector(to_unsigned(1328, LDPC_TABLE_DATA_WIDTH)),
    6440 => std_logic_vector(to_unsigned(329, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6441 => std_logic_vector(to_unsigned(3, LDPC_TABLE_DATA_WIDTH)),
    6442 => std_logic_vector(to_unsigned(1515, LDPC_TABLE_DATA_WIDTH)),
    6443 => std_logic_vector(to_unsigned(506, LDPC_TABLE_DATA_WIDTH)), -- last item of row
    6444 => std_logic_vector(to_unsigned(4, LDPC_TABLE_DATA_WIDTH)),
    6445 => std_logic_vector(to_unsigned(1104, LDPC_TABLE_DATA_WIDTH)),
    6446 => std_logic_vector(to_unsigned(1172, LDPC_TABLE_DATA_WIDTH)));

end package ldpc_tables_pkg;

package body ldpc_tables_pkg is
  -- Use this function to get the starting address of a given config within the LDPC_DATA_TABLE
  function get_ldpc_metadata (
    constant frame_length : frame_type_t;
    constant code_rate : code_rate_t) return ldpc_metadata_t is
  begin
    if frame_length = fecframe_normal and code_rate = C1_2 then
      return (
        addr => 0,
        q => 90,
        stage_0_loops => 36,
        stage_0_rows => 8,
        stage_1_loops => 54,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C1_3 then
      return (
        addr => 450,
        q => 120,
        stage_0_loops => 20,
        stage_0_rows => 12,
        stage_1_loops => 40,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C1_4 then
      return (
        addr => 810,
        q => 135,
        stage_0_loops => 15,
        stage_0_rows => 12,
        stage_1_loops => 30,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C2_3 then
      return (
        addr => 1080,
        q => 60,
        stage_0_loops => 12,
        stage_0_rows => 13,
        stage_1_loops => 108,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C2_5 then
      return (
        addr => 1560,
        q => 108,
        stage_0_loops => 24,
        stage_0_rows => 12,
        stage_1_loops => 48,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C3_4 then
      return (
        addr => 1992,
        q => 45,
        stage_0_loops => 15,
        stage_0_rows => 12,
        stage_1_loops => 120,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C3_5 then
      return (
        addr => 2532,
        q => 72,
        stage_0_loops => 36,
        stage_0_rows => 12,
        stage_1_loops => 72,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C4_5 then
      return (
        addr => 3180,
        q => 36,
        stage_0_loops => 18,
        stage_0_rows => 11,
        stage_1_loops => 126,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C5_6 then
      return (
        addr => 3756,
        q => 30,
        stage_0_loops => 15,
        stage_0_rows => 13,
        stage_1_loops => 135,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C8_9 then
      return (
        addr => 4356,
        q => 20,
        stage_0_loops => 20,
        stage_0_rows => 4,
        stage_1_loops => 140,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_normal and code_rate = C9_10 then
      return (
        addr => 4856,
        q => 18,
        stage_0_loops => 18,
        stage_0_rows => 4,
        stage_1_loops => 144,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_2 then
      return (
        addr => 5360,
        q => 25,
        stage_0_loops => 5,
        stage_0_rows => 8,
        stage_1_loops => 15,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_3 then
      return (
        addr => 5445,
        q => 30,
        stage_0_loops => 5,
        stage_0_rows => 12,
        stage_1_loops => 10,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C1_4 then
      return (
        addr => 5535,
        q => 36,
        stage_0_loops => 4,
        stage_0_rows => 12,
        stage_1_loops => 5,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C2_3 then
      return (
        addr => 5598,
        q => 15,
        stage_0_loops => 3,
        stage_0_rows => 13,
        stage_1_loops => 27,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C2_5 then
      return (
        addr => 5718,
        q => 27,
        stage_0_loops => 6,
        stage_0_rows => 12,
        stage_1_loops => 12,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C3_4 then
      return (
        addr => 5826,
        q => 12,
        stage_0_loops => 1,
        stage_0_rows => 12,
        stage_1_loops => 32,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C3_5 then
      return (
        addr => 5934,
        q => 18,
        stage_0_loops => 9,
        stage_0_rows => 12,
        stage_1_loops => 18,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C4_5 then
      return (
        addr => 6096,
        q => 10,
        stage_0_loops => 17,
        stage_0_rows => 3,
        stage_1_loops => 18,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C5_6 then
      return (
        addr => 6201,
        q => 8,
        stage_0_loops => 1,
        stage_0_rows => 13,
        stage_1_loops => 36,
        stage_1_rows => 3);
     end if;
    if frame_length = fecframe_short and code_rate = C8_9 then
      return (
        addr => 6322,
        q => 5,
        stage_0_loops => 5,
        stage_0_rows => 4,
        stage_1_loops => 35,
        stage_1_rows => 3);
     end if;

    -- Return a non existing index for any config not listed above
    return (addr => -1, q => -1, stage_0_loops => -1, stage_0_rows => -1, stage_1_loops => -1, stage_1_rows => -1);
  end function get_ldpc_metadata;

end package body ldpc_tables_pkg;