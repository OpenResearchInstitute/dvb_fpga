--
-- DVB IP
--
-- Copyright 2020 by Suoto <andre820@gmail.com>
--
-- This file is part of the DVB IP.
--
-- DVB IP is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- DVB IP is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with DVB IP.  If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library fpga_cores;
use fpga_cores.common_pkg.all;

-- Summary of statistics

--    table                               depth    width (bits)    width (entries)    total (bytes)    18k BRAMs    36k BRAMs
----  --------------------------------  -------  --------------  -----------------  ---------------  -----------  -----------
--    ldpc_table_FECFRAME_NORMAL_C1_2        90             115                  9             1294            7            4
--    ldpc_table_FECFRAME_NORMAL_C1_3        60             196                 13             1470           11            6
--    ldpc_table_FECFRAME_NORMAL_C1_4        45             196                 13             1103           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_3       120             189                 14             2835           11            6
--    ldpc_table_FECFRAME_NORMAL_C2_5        72             196                 13             1764           11            6
--    ldpc_table_FECFRAME_NORMAL_C3_4       135             164                 13             2768           10            5
--    ldpc_table_FECFRAME_NORMAL_C3_5       108             184                 13             2484           11            6
--    ldpc_table_FECFRAME_NORMAL_C4_5       144             150                 12             2700            9            5
--    ldpc_table_FECFRAME_NORMAL_C5_6       150             177                 14             3319           10            5
--    ldpc_table_FECFRAME_NORMAL_C8_9       160              46                  5              920            3            2
--    ldpc_table_FECFRAME_NORMAL_C9_10      162              46                  5              932            3            2
--    ldpc_table_FECFRAME_SHORT_C1_2         20             100                  9              250            6            3
--    ldpc_table_FECFRAME_SHORT_C1_3         15             170                 13              319           10            5
--    ldpc_table_FECFRAME_SHORT_C1_4          9             171                 13              193           10            5
--    ldpc_table_FECFRAME_SHORT_C2_3         30             156                 14              585            9            5
--    ldpc_table_FECFRAME_SHORT_C2_5         18             168                 13              378           10            5
--    ldpc_table_FECFRAME_SHORT_C3_4         33             133                 13              549            8            4
--    ldpc_table_FECFRAME_SHORT_C3_5         27             160                 13              540            9            5
--    ldpc_table_FECFRAME_SHORT_C4_5         35              30                  4              132            2            1
--    ldpc_table_FECFRAME_SHORT_C5_6         37             139                 14              643            8            4
--    ldpc_table_FECFRAME_SHORT_C8_9         40              37                  5              185            3            2

package ldpc_tables_pkg is

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_2.csv, table is 90x115 (1293.75 bytes)
  -- Resource estimation: 7 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 7, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_2 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 89)(0 to 8)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 8, 1 => 54, 2 => 9318, 3 => 14392, 4 => 27561, 5 => 26909, 6 => 10219, 7 => 2534, 8 => 8597),
    1 => integer_vector_t'(0 => 8, 1 => 55, 2 => 7263, 3 => 4635, 4 => 2530, 5 => 28130, 6 => 3033, 7 => 23830, 8 => 3651),
    2 => integer_vector_t'(0 => 8, 1 => 56, 2 => 24731, 3 => 23583, 4 => 26036, 5 => 17299, 6 => 5750, 7 => 792, 8 => 9169),
    3 => integer_vector_t'(0 => 8, 1 => 57, 2 => 5811, 3 => 26154, 4 => 18653, 5 => 11551, 6 => 15447, 7 => 13685, 8 => 16264),
    4 => integer_vector_t'(0 => 8, 1 => 58, 2 => 12610, 3 => 11347, 4 => 28768, 5 => 2792, 6 => 3174, 7 => 29371, 8 => 12997),
    5 => integer_vector_t'(0 => 8, 1 => 59, 2 => 16789, 3 => 16018, 4 => 21449, 5 => 6165, 6 => 21202, 7 => 15850, 8 => 3186),
    6 => integer_vector_t'(0 => 8, 1 => 60, 2 => 31016, 3 => 21449, 4 => 17618, 5 => 6213, 6 => 12166, 7 => 8334, 8 => 18212),
    7 => integer_vector_t'(0 => 8, 1 => 61, 2 => 22836, 3 => 14213, 4 => 11327, 5 => 5896, 6 => 718, 7 => 11727, 8 => 9308),
    8 => integer_vector_t'(0 => 8, 1 => 62, 2 => 2091, 3 => 24941, 4 => 29966, 5 => 23634, 6 => 9013, 7 => 15587, 8 => 5444),
    9 => integer_vector_t'(0 => 8, 1 => 63, 2 => 22207, 3 => 3983, 4 => 16904, 5 => 28534, 6 => 21415, 7 => 27524, 8 => 25912),
    10 => integer_vector_t'(0 => 8, 1 => 64, 2 => 25687, 3 => 4501, 4 => 22193, 5 => 14665, 6 => 14798, 7 => 16158, 8 => 5491),
    11 => integer_vector_t'(0 => 8, 1 => 65, 2 => 4520, 3 => 17094, 4 => 23397, 5 => 4264, 6 => 22370, 7 => 16941, 8 => 21526),
    12 => integer_vector_t'(0 => 8, 1 => 66, 2 => 10490, 3 => 6182, 4 => 32370, 5 => 9597, 6 => 30841, 7 => 25954, 8 => 2762),
    13 => integer_vector_t'(0 => 8, 1 => 67, 2 => 22120, 3 => 22865, 4 => 29870, 5 => 15147, 6 => 13668, 7 => 14955, 8 => 19235),
    14 => integer_vector_t'(0 => 8, 1 => 68, 2 => 6689, 3 => 18408, 4 => 18346, 5 => 9918, 6 => 25746, 7 => 5443, 8 => 20645),
    15 => integer_vector_t'(0 => 8, 1 => 69, 2 => 29982, 3 => 12529, 4 => 13858, 5 => 4746, 6 => 30370, 7 => 10023, 8 => 24828),
    16 => integer_vector_t'(0 => 8, 1 => 70, 2 => 1262, 3 => 28032, 4 => 29888, 5 => 13063, 6 => 24033, 7 => 21951, 8 => 7863),
    17 => integer_vector_t'(0 => 8, 1 => 71, 2 => 6594, 3 => 29642, 4 => 31451, 5 => 14831, 6 => 9509, 7 => 9335, 8 => 31552),
    18 => integer_vector_t'(0 => 8, 1 => 72, 2 => 1358, 3 => 6454, 4 => 16633, 5 => 20354, 6 => 24598, 7 => 624, 8 => 5265),
    19 => integer_vector_t'(0 => 8, 1 => 73, 2 => 19529, 3 => 295, 4 => 18011, 5 => 3080, 6 => 13364, 7 => 8032, 8 => 15323),
    20 => integer_vector_t'(0 => 8, 1 => 74, 2 => 11981, 3 => 1510, 4 => 7960, 5 => 21462, 6 => 9129, 7 => 11370, 8 => 25741),
    21 => integer_vector_t'(0 => 8, 1 => 75, 2 => 9276, 3 => 29656, 4 => 4543, 5 => 30699, 6 => 20646, 7 => 21921, 8 => 28050),
    22 => integer_vector_t'(0 => 8, 1 => 76, 2 => 15975, 3 => 25634, 4 => 5520, 5 => 31119, 6 => 13715, 7 => 21949, 8 => 19605),
    23 => integer_vector_t'(0 => 8, 1 => 77, 2 => 18688, 3 => 4608, 4 => 31755, 5 => 30165, 6 => 13103, 7 => 10706, 8 => 29224),
    24 => integer_vector_t'(0 => 8, 1 => 78, 2 => 21514, 3 => 23117, 4 => 12245, 5 => 26035, 6 => 31656, 7 => 25631, 8 => 30699),
    25 => integer_vector_t'(0 => 8, 1 => 79, 2 => 9674, 3 => 24966, 4 => 31285, 5 => 29908, 6 => 17042, 7 => 24588, 8 => 31857),
    26 => integer_vector_t'(0 => 8, 1 => 80, 2 => 21856, 3 => 27777, 4 => 29919, 5 => 27000, 6 => 14897, 7 => 11409, 8 => 7122),
    27 => integer_vector_t'(0 => 8, 1 => 81, 2 => 29773, 3 => 23310, 4 => 263, 5 => 4877, 6 => 28622, 7 => 20545, 8 => 22092),
    28 => integer_vector_t'(0 => 8, 1 => 82, 2 => 15605, 3 => 5651, 4 => 21864, 5 => 3967, 6 => 14419, 7 => 22757, 8 => 15896),
    29 => integer_vector_t'(0 => 8, 1 => 83, 2 => 30145, 3 => 1759, 4 => 10139, 5 => 29223, 6 => 26086, 7 => 10556, 8 => 5098),
    30 => integer_vector_t'(0 => 8, 1 => 84, 2 => 18815, 3 => 16575, 4 => 2936, 5 => 24457, 6 => 26738, 7 => 6030, 8 => 505),
    31 => integer_vector_t'(0 => 8, 1 => 85, 2 => 30326, 3 => 22298, 4 => 27562, 5 => 20131, 6 => 26390, 7 => 6247, 8 => 24791),
    32 => integer_vector_t'(0 => 8, 1 => 86, 2 => 928, 3 => 29246, 4 => 21246, 5 => 12400, 6 => 15311, 7 => 32309, 8 => 18608),
    33 => integer_vector_t'(0 => 8, 1 => 87, 2 => 20314, 3 => 6025, 4 => 26689, 5 => 16302, 6 => 2296, 7 => 3244, 8 => 19613),
    34 => integer_vector_t'(0 => 8, 1 => 88, 2 => 6237, 3 => 11943, 4 => 22851, 5 => 15642, 6 => 23857, 7 => 15112, 8 => 20947),
    35 => integer_vector_t'(0 => 8, 1 => 89, 2 => 26403, 3 => 25168, 4 => 19038, 5 => 18384, 6 => 8882, 7 => 12719, 8 => 7093),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 14567, 3 => 24965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3908, 3 => 100, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10279, 3 => 240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 24102, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 12383, 3 => 4173, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 13861, 3 => 15918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 21327, 3 => 1046, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5288, 3 => 14579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 28158, 3 => 8069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 16583, 3 => 11098, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 16681, 3 => 28363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 13980, 3 => 24725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 32169, 3 => 17989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 10907, 3 => 2767, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 21557, 3 => 3818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 26676, 3 => 12422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 7676, 3 => 8754, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 14905, 3 => 20232, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 15719, 3 => 24646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 31942, 3 => 8589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 19978, 3 => 27197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 27060, 3 => 15071, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6071, 3 => 26649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10393, 3 => 11176, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 9597, 3 => 13370, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7081, 3 => 17677, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 1433, 3 => 19513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 26925, 3 => 9014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 19202, 3 => 8900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 18152, 3 => 30647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20803, 3 => 1737, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 11804, 3 => 25221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 31683, 3 => 17783, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 29694, 3 => 9345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 12280, 3 => 26611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 6526, 3 => 26122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 26165, 3 => 11241, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 7666, 3 => 26962, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 16290, 3 => 8480, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 11774, 3 => 10120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 30051, 3 => 30426, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 1335, 3 => 15424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6865, 3 => 17742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 31779, 3 => 12489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 32120, 3 => 21001, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 14508, 3 => 6996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 979, 3 => 25024, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 4554, 3 => 21896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 7989, 3 => 21777, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 4972, 3 => 20661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 6612, 3 => 2730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 12742, 3 => 4418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 29194, 3 => 595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 19267, 3 => 20113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_3.csv, table is 60x196 (1470.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_3 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 59)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 34903, 2 => 20927, 3 => 32093, 4 => 1052, 5 => 25611, 6 => 16093, 7 => 16454, 8 => 5520, 9 => 506, 10 => 37399, 11 => 18518, 12 => 21120),
    1 => integer_vector_t'(0 => 12, 1 => 11636, 2 => 14594, 3 => 22158, 4 => 14763, 5 => 15333, 6 => 6838, 7 => 22222, 8 => 37856, 9 => 14985, 10 => 31041, 11 => 18704, 12 => 32910),
    2 => integer_vector_t'(0 => 12, 1 => 17449, 2 => 1665, 3 => 35639, 4 => 16624, 5 => 12867, 6 => 12449, 7 => 10241, 8 => 11650, 9 => 25622, 10 => 34372, 11 => 19878, 12 => 26894),
    3 => integer_vector_t'(0 => 12, 1 => 29235, 2 => 19780, 3 => 36056, 4 => 20129, 5 => 20029, 6 => 5457, 7 => 8157, 8 => 35554, 9 => 21237, 10 => 7943, 11 => 13873, 12 => 14980),
    4 => integer_vector_t'(0 => 12, 1 => 9912, 2 => 7143, 3 => 35911, 4 => 12043, 5 => 17360, 6 => 37253, 7 => 25588, 8 => 11827, 9 => 29152, 10 => 21936, 11 => 24125, 12 => 40870),
    5 => integer_vector_t'(0 => 12, 1 => 40701, 2 => 36035, 3 => 39556, 4 => 12366, 5 => 19946, 6 => 29072, 7 => 16365, 8 => 35495, 9 => 22686, 10 => 11106, 11 => 8756, 12 => 34863),
    6 => integer_vector_t'(0 => 12, 1 => 19165, 2 => 15702, 3 => 13536, 4 => 40238, 5 => 4465, 6 => 40034, 7 => 40590, 8 => 37540, 9 => 17162, 10 => 1712, 11 => 20577, 12 => 14138),
    7 => integer_vector_t'(0 => 12, 1 => 31338, 2 => 19342, 3 => 9301, 4 => 39375, 5 => 3211, 6 => 1316, 7 => 33409, 8 => 28670, 9 => 12282, 10 => 6118, 11 => 29236, 12 => 35787),
    8 => integer_vector_t'(0 => 12, 1 => 11504, 2 => 30506, 3 => 19558, 4 => 5100, 5 => 24188, 6 => 24738, 7 => 30397, 8 => 33775, 9 => 9699, 10 => 6215, 11 => 3397, 12 => 37451),
    9 => integer_vector_t'(0 => 12, 1 => 34689, 2 => 23126, 3 => 7571, 4 => 1058, 5 => 12127, 6 => 27518, 7 => 23064, 8 => 11265, 9 => 14867, 10 => 30451, 11 => 28289, 12 => 2966),
    10 => integer_vector_t'(0 => 12, 1 => 11660, 2 => 15334, 3 => 16867, 4 => 15160, 5 => 38343, 6 => 3778, 7 => 4265, 8 => 39139, 9 => 17293, 10 => 26229, 11 => 42604, 12 => 13486),
    11 => integer_vector_t'(0 => 12, 1 => 31497, 2 => 1365, 3 => 14828, 4 => 7453, 5 => 26350, 6 => 41346, 7 => 28643, 8 => 23421, 9 => 8354, 10 => 16255, 11 => 11055, 12 => 24279),
    12 => integer_vector_t'(0 => 12, 1 => 15687, 2 => 12467, 3 => 13906, 4 => 5215, 5 => 41328, 6 => 23755, 7 => 20800, 8 => 6447, 9 => 7970, 10 => 2803, 11 => 33262, 12 => 39843),
    13 => integer_vector_t'(0 => 12, 1 => 5363, 2 => 22469, 3 => 38091, 4 => 28457, 5 => 36696, 6 => 34471, 7 => 23619, 8 => 2404, 9 => 24229, 10 => 41754, 11 => 1297, 12 => 18563),
    14 => integer_vector_t'(0 => 12, 1 => 3673, 2 => 39070, 3 => 14480, 4 => 30279, 5 => 37483, 6 => 7580, 7 => 29519, 8 => 30519, 9 => 39831, 10 => 20252, 11 => 18132, 12 => 20010),
    15 => integer_vector_t'(0 => 12, 1 => 34386, 2 => 7252, 3 => 27526, 4 => 12950, 5 => 6875, 6 => 43020, 7 => 31566, 8 => 39069, 9 => 18985, 10 => 15541, 11 => 40020, 12 => 16715),
    16 => integer_vector_t'(0 => 12, 1 => 1721, 2 => 37332, 3 => 39953, 4 => 17430, 5 => 32134, 6 => 29162, 7 => 10490, 8 => 12971, 9 => 28581, 10 => 29331, 11 => 6489, 12 => 35383),
    17 => integer_vector_t'(0 => 12, 1 => 736, 2 => 7022, 3 => 42349, 4 => 8783, 5 => 6767, 6 => 11871, 7 => 21675, 8 => 10325, 9 => 11548, 10 => 25978, 11 => 431, 12 => 24085),
    18 => integer_vector_t'(0 => 12, 1 => 1925, 2 => 10602, 3 => 28585, 4 => 12170, 5 => 15156, 6 => 34404, 7 => 8351, 8 => 13273, 9 => 20208, 10 => 5800, 11 => 15367, 12 => 21764),
    19 => integer_vector_t'(0 => 12, 1 => 16279, 2 => 37832, 3 => 34792, 4 => 21250, 5 => 34192, 6 => 7406, 7 => 41488, 8 => 18346, 9 => 29227, 10 => 26127, 11 => 25493, 12 => 7048),
    20 => integer_vector_t'(0 => 3, 1 => 39948, 2 => 28229, 3 => 24899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 17408, 2 => 14274, 3 => 38993, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 38774, 2 => 15968, 3 => 28459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 41404, 2 => 27249, 3 => 27425, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 41229, 2 => 6082, 3 => 43114, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 13957, 2 => 4979, 3 => 40654, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 3093, 2 => 3438, 3 => 34992, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 34082, 2 => 6172, 3 => 28760, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 42210, 2 => 34141, 3 => 41021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14705, 2 => 17783, 3 => 10134, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 41755, 2 => 39884, 3 => 22773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14615, 2 => 15593, 3 => 1642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 29111, 2 => 37061, 3 => 39860, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 9579, 2 => 33552, 3 => 633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 12951, 2 => 21137, 3 => 39608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 38244, 2 => 27361, 3 => 29417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 2939, 2 => 10172, 3 => 36479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 29094, 2 => 5357, 3 => 19224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 9562, 2 => 24436, 3 => 28637, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 40177, 2 => 2326, 3 => 13504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 6834, 2 => 21583, 3 => 42516, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 40651, 2 => 42810, 3 => 25709, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 31557, 2 => 32138, 3 => 38142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 18624, 2 => 41867, 3 => 39296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 37560, 2 => 14295, 3 => 16245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 6821, 2 => 21679, 3 => 31570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 25339, 2 => 25083, 3 => 22081, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 8047, 2 => 697, 3 => 35268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 9884, 2 => 17073, 3 => 19995, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 26848, 2 => 35245, 3 => 8390, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 18658, 2 => 16134, 3 => 14807, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 12201, 2 => 32944, 3 => 5035, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 25236, 2 => 1216, 3 => 38986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 42994, 2 => 24782, 3 => 8681, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 28321, 2 => 4932, 3 => 34249, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 4107, 2 => 29382, 3 => 32124, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 22157, 2 => 2624, 3 => 14468, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 38788, 2 => 27081, 3 => 7936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4368, 2 => 26148, 3 => 10578, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 25353, 2 => 4122, 3 => 39751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C1_4.csv, table is 45x196 (1102.5 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C1_4 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 44)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 23606, 2 => 36098, 3 => 1140, 4 => 28859, 5 => 18148, 6 => 18510, 7 => 6226, 8 => 540, 9 => 42014, 10 => 20879, 11 => 23802, 12 => 47088),
    1 => integer_vector_t'(0 => 12, 1 => 16419, 2 => 24928, 3 => 16609, 4 => 17248, 5 => 7693, 6 => 24997, 7 => 42587, 8 => 16858, 9 => 34921, 10 => 21042, 11 => 37024, 12 => 20692),
    2 => integer_vector_t'(0 => 12, 1 => 1874, 2 => 40094, 3 => 18704, 4 => 14474, 5 => 14004, 6 => 11519, 7 => 13106, 8 => 28826, 9 => 38669, 10 => 22363, 11 => 30255, 12 => 31105),
    3 => integer_vector_t'(0 => 12, 1 => 22254, 2 => 40564, 3 => 22645, 4 => 22532, 5 => 6134, 6 => 9176, 7 => 39998, 8 => 23892, 9 => 8937, 10 => 15608, 11 => 16854, 12 => 31009),
    4 => integer_vector_t'(0 => 12, 1 => 8037, 2 => 40401, 3 => 13550, 4 => 19526, 5 => 41902, 6 => 28782, 7 => 13304, 8 => 32796, 9 => 24679, 10 => 27140, 11 => 45980, 12 => 10021),
    5 => integer_vector_t'(0 => 12, 1 => 40540, 2 => 44498, 3 => 13911, 4 => 22435, 5 => 32701, 6 => 18405, 7 => 39929, 8 => 25521, 9 => 12497, 10 => 9851, 11 => 39223, 12 => 34823),
    6 => integer_vector_t'(0 => 12, 1 => 15233, 2 => 45333, 3 => 5041, 4 => 44979, 5 => 45710, 6 => 42150, 7 => 19416, 8 => 1892, 9 => 23121, 10 => 15860, 11 => 8832, 12 => 10308),
    7 => integer_vector_t'(0 => 12, 1 => 10468, 2 => 44296, 3 => 3611, 4 => 1480, 5 => 37581, 6 => 32254, 7 => 13817, 8 => 6883, 9 => 32892, 10 => 40258, 11 => 46538, 12 => 11940),
    8 => integer_vector_t'(0 => 12, 1 => 6705, 2 => 21634, 3 => 28150, 4 => 43757, 5 => 895, 6 => 6547, 7 => 20970, 8 => 28914, 9 => 30117, 10 => 25736, 11 => 41734, 12 => 11392),
    9 => integer_vector_t'(0 => 12, 1 => 22002, 2 => 5739, 3 => 27210, 4 => 27828, 5 => 34192, 6 => 37992, 7 => 10915, 8 => 6998, 9 => 3824, 10 => 42130, 11 => 4494, 12 => 35739),
    10 => integer_vector_t'(0 => 12, 1 => 8515, 2 => 1191, 3 => 13642, 4 => 30950, 5 => 25943, 6 => 12673, 7 => 16726, 8 => 34261, 9 => 31828, 10 => 3340, 11 => 8747, 12 => 39225),
    11 => integer_vector_t'(0 => 12, 1 => 18979, 2 => 17058, 3 => 43130, 4 => 4246, 5 => 4793, 6 => 44030, 7 => 19454, 8 => 29511, 9 => 47929, 10 => 15174, 11 => 24333, 12 => 19354),
    12 => integer_vector_t'(0 => 12, 1 => 16694, 2 => 8381, 3 => 29642, 4 => 46516, 5 => 32224, 6 => 26344, 7 => 9405, 8 => 18292, 9 => 12437, 10 => 27316, 11 => 35466, 12 => 41992),
    13 => integer_vector_t'(0 => 12, 1 => 15642, 2 => 5871, 3 => 46489, 4 => 26723, 5 => 23396, 6 => 7257, 7 => 8974, 8 => 3156, 9 => 37420, 10 => 44823, 11 => 35423, 12 => 13541),
    14 => integer_vector_t'(0 => 12, 1 => 42858, 2 => 32008, 3 => 41282, 4 => 38773, 5 => 26570, 6 => 2702, 7 => 27260, 8 => 46974, 9 => 1469, 10 => 20887, 11 => 27426, 12 => 38553),
    15 => integer_vector_t'(0 => 3, 1 => 22152, 2 => 24261, 3 => 8297, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 19347, 2 => 9978, 3 => 27802, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 34991, 2 => 6354, 3 => 33561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 29782, 2 => 30875, 3 => 29523, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 9278, 2 => 48512, 3 => 14349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 38061, 2 => 4165, 3 => 43878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 8548, 2 => 33172, 3 => 34410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22535, 2 => 28811, 3 => 23950, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 20439, 2 => 4027, 3 => 24186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 38618, 2 => 8187, 3 => 30947, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 35538, 2 => 43880, 3 => 21459, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 7091, 2 => 45616, 3 => 15063, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 5505, 2 => 9315, 3 => 21908, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 36046, 2 => 32914, 3 => 11836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 7304, 2 => 39782, 3 => 33721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 16905, 2 => 29962, 3 => 12980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11171, 2 => 23709, 3 => 22460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 34541, 2 => 9937, 3 => 44500, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 14035, 2 => 47316, 3 => 8815, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 15057, 2 => 45482, 3 => 24461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 30518, 2 => 36877, 3 => 879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7583, 2 => 13364, 3 => 24332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 448, 2 => 27056, 3 => 4682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 12083, 2 => 31378, 3 => 21670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 1159, 2 => 18031, 3 => 2221, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 17028, 2 => 38715, 3 => 9350, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 17343, 2 => 24530, 3 => 29574, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 46128, 2 => 31039, 3 => 32818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 20373, 2 => 36967, 3 => 18345, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 46685, 2 => 20622, 3 => 32806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_3.csv, table is 120x189 (2835.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 14, 9 => 15, 10 => 15, 11 => 15, 12 => 15, 13 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_3 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 119)(0 to 13)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 10491, 3 => 16043, 4 => 506, 5 => 12826, 6 => 8065, 7 => 8226, 8 => 2767, 9 => 240, 10 => 18673, 11 => 9279, 12 => 10579, 13 => 20928),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 17819, 3 => 8313, 4 => 6433, 5 => 6224, 6 => 5120, 7 => 5824, 8 => 12812, 9 => 17187, 10 => 9940, 11 => 13447, 12 => 13825, 13 => 18483),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 17957, 3 => 6024, 4 => 8681, 5 => 18628, 6 => 12794, 7 => 5915, 8 => 14576, 9 => 10970, 10 => 12064, 11 => 20437, 12 => 4455, 13 => 7151),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 19777, 3 => 6183, 4 => 9972, 5 => 14536, 6 => 8182, 7 => 17749, 8 => 11341, 9 => 5556, 10 => 4379, 11 => 17434, 12 => 15477, 13 => 18532),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 4651, 3 => 19689, 4 => 1608, 5 => 659, 6 => 16707, 7 => 14335, 8 => 6143, 9 => 3058, 10 => 14618, 11 => 17894, 12 => 20684, 13 => 5306),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 9778, 3 => 2552, 4 => 12096, 5 => 12369, 6 => 15198, 7 => 16890, 8 => 4851, 9 => 3109, 10 => 1700, 11 => 18725, 12 => 1997, 13 => 15882),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 486, 3 => 6111, 4 => 13743, 5 => 11537, 6 => 5591, 7 => 7433, 8 => 15227, 9 => 14145, 10 => 1483, 11 => 3887, 12 => 17431, 13 => 12430),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 20647, 3 => 14311, 4 => 11734, 5 => 4180, 6 => 8110, 7 => 5525, 8 => 12141, 9 => 15761, 10 => 18661, 11 => 18441, 12 => 10569, 13 => 8192),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 3791, 3 => 14759, 4 => 15264, 5 => 19918, 6 => 10132, 7 => 9062, 8 => 10010, 9 => 12786, 10 => 10675, 11 => 9682, 12 => 19246, 13 => 5454),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 19525, 3 => 9485, 4 => 7777, 5 => 19999, 6 => 8378, 7 => 9209, 8 => 3163, 9 => 20232, 10 => 6690, 11 => 16518, 12 => 716, 13 => 7353),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 4588, 3 => 6709, 4 => 20202, 5 => 10905, 6 => 915, 7 => 4317, 8 => 11073, 9 => 13576, 10 => 16433, 11 => 368, 12 => 3508, 13 => 21171),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 14072, 3 => 4033, 4 => 19959, 5 => 12608, 6 => 631, 7 => 19494, 8 => 14160, 9 => 8249, 10 => 10223, 11 => 21504, 12 => 12395, 13 => 4322),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 13800, 3 => 14161, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2948, 3 => 9647, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 14693, 3 => 16027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 20506, 3 => 11082, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1143, 3 => 9020, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13501, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1548, 3 => 2190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 12216, 3 => 21556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 19897, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4189, 3 => 7958, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 15940, 3 => 10048, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 515, 3 => 12614, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8501, 3 => 8450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 17595, 3 => 16784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 5913, 3 => 8495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 16394, 3 => 10423, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7409, 3 => 6981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6678, 3 => 15939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 20344, 3 => 12987, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 2510, 3 => 14588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 17918, 3 => 6655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 6703, 3 => 19451, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 496, 3 => 4217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7290, 3 => 5766, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 10521, 3 => 8925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 20379, 3 => 11905, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4090, 3 => 5838, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 19082, 3 => 17040, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 20233, 3 => 12352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 19365, 3 => 19546, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 6249, 3 => 19030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11037, 3 => 19193, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 19760, 3 => 11772, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 45, 2 => 19644, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16076, 3 => 3521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11779, 3 => 21062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 48, 2 => 13062, 3 => 9682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 49, 2 => 8934, 3 => 5217, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 50, 2 => 11087, 3 => 3319, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 51, 2 => 18892, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 52, 2 => 7894, 3 => 3898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 53, 2 => 5963, 3 => 4360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 54, 2 => 7346, 3 => 11726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5182, 3 => 5609, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 56, 2 => 2412, 3 => 17295, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 57, 2 => 9845, 3 => 20494, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 58, 2 => 6687, 3 => 1864, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 59, 2 => 20564, 3 => 5216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18226, 3 => 17207, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9380, 3 => 8266, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7073, 3 => 3065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 18252, 3 => 13437, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9161, 3 => 15642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10714, 3 => 10153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 11585, 3 => 9078, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5359, 3 => 9418, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 9024, 3 => 9515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1206, 3 => 16354, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 14994, 3 => 1102, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9375, 3 => 20796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 15964, 3 => 6027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14789, 3 => 6452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8002, 3 => 18591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 14742, 3 => 14089, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 253, 3 => 3045, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1274, 3 => 19286, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 14777, 3 => 2044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 13920, 3 => 9900, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 452, 3 => 7374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 18206, 3 => 9921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6131, 3 => 5414, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10077, 3 => 9726, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 12045, 3 => 5479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4322, 3 => 7990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 15616, 3 => 5550, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 15561, 3 => 10661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 20718, 3 => 7387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2518, 3 => 18804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8984, 3 => 2600, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6516, 3 => 17909, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 32, 2 => 11148, 3 => 98, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 33, 2 => 20559, 3 => 3704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7510, 3 => 1569, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 35, 2 => 16000, 3 => 11692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 36, 2 => 9147, 3 => 10303, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 37, 2 => 16650, 3 => 191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15577, 3 => 18685, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 39, 2 => 17167, 3 => 20917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 40, 2 => 4256, 3 => 3391, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 41, 2 => 20092, 3 => 17219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 42, 2 => 9218, 3 => 5056, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 43, 2 => 18429, 3 => 8472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12093, 3 => 20753, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 45, 2 => 16345, 3 => 12748, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 46, 2 => 16023, 3 => 11095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 47, 2 => 5048, 3 => 17595, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 48, 2 => 18995, 3 => 4817, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 49, 2 => 16483, 3 => 3536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 50, 2 => 1439, 3 => 16148, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 51, 2 => 3661, 3 => 3039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 52, 2 => 19010, 3 => 18121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 53, 2 => 8968, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 54, 2 => 13427, 3 => 18003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 55, 2 => 5303, 3 => 3083, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 56, 2 => 531, 3 => 16668, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 57, 2 => 4771, 3 => 6722, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 58, 2 => 5695, 3 => 7960, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 59, 2 => 3589, 3 => 14630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C2_5.csv, table is 72x196 (1764.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant LDPC_TABLE_FECFRAME_NORMAL_C2_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 71)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 31413, 2 => 18834, 3 => 28884, 4 => 947, 5 => 23050, 6 => 14484, 7 => 14809, 8 => 4968, 9 => 455, 10 => 33659, 11 => 16666, 12 => 19008),
    1 => integer_vector_t'(0 => 12, 1 => 13172, 2 => 19939, 3 => 13354, 4 => 13719, 5 => 6132, 6 => 20086, 7 => 34040, 8 => 13442, 9 => 27958, 10 => 16813, 11 => 29619, 12 => 16553),
    2 => integer_vector_t'(0 => 12, 1 => 1499, 2 => 32075, 3 => 14962, 4 => 11578, 5 => 11204, 6 => 9217, 7 => 10485, 8 => 23062, 9 => 30936, 10 => 17892, 11 => 24204, 12 => 24885),
    3 => integer_vector_t'(0 => 12, 1 => 32490, 2 => 18086, 3 => 18007, 4 => 4957, 5 => 7285, 6 => 32073, 7 => 19038, 8 => 7152, 9 => 12486, 10 => 13483, 11 => 24808, 12 => 21759),
    4 => integer_vector_t'(0 => 12, 1 => 32321, 2 => 10839, 3 => 15620, 4 => 33521, 5 => 23030, 6 => 10646, 7 => 26236, 8 => 19744, 9 => 21713, 10 => 36784, 11 => 8016, 12 => 12869),
    5 => integer_vector_t'(0 => 12, 1 => 35597, 2 => 11129, 3 => 17948, 4 => 26160, 5 => 14729, 6 => 31943, 7 => 20416, 8 => 10000, 9 => 7882, 10 => 31380, 11 => 27858, 12 => 33356),
    6 => integer_vector_t'(0 => 12, 1 => 14125, 2 => 12131, 3 => 36199, 4 => 4058, 5 => 35992, 6 => 36594, 7 => 33698, 8 => 15475, 9 => 1566, 10 => 18498, 11 => 12725, 12 => 7067),
    7 => integer_vector_t'(0 => 12, 1 => 17406, 2 => 8372, 3 => 35437, 4 => 2888, 5 => 1184, 6 => 30068, 7 => 25802, 8 => 11056, 9 => 5507, 10 => 26313, 11 => 32205, 12 => 37232),
    8 => integer_vector_t'(0 => 12, 1 => 15254, 2 => 5365, 3 => 17308, 4 => 22519, 5 => 35009, 6 => 718, 7 => 5240, 8 => 16778, 9 => 23131, 10 => 24092, 11 => 20587, 12 => 33385),
    9 => integer_vector_t'(0 => 12, 1 => 27455, 2 => 17602, 3 => 4590, 4 => 21767, 5 => 22266, 6 => 27357, 7 => 30400, 8 => 8732, 9 => 5596, 10 => 3060, 11 => 33703, 12 => 3596),
    10 => integer_vector_t'(0 => 12, 1 => 6882, 2 => 873, 3 => 10997, 4 => 24738, 5 => 20770, 6 => 10067, 7 => 13379, 8 => 27409, 9 => 25463, 10 => 2673, 11 => 6998, 12 => 31378),
    11 => integer_vector_t'(0 => 12, 1 => 15181, 2 => 13645, 3 => 34501, 4 => 3393, 5 => 3840, 6 => 35227, 7 => 15562, 8 => 23615, 9 => 38342, 10 => 12139, 11 => 19471, 12 => 15483),
    12 => integer_vector_t'(0 => 12, 1 => 13350, 2 => 6707, 3 => 23709, 4 => 37204, 5 => 25778, 6 => 21082, 7 => 7511, 8 => 14588, 9 => 10010, 10 => 21854, 11 => 28375, 12 => 33591),
    13 => integer_vector_t'(0 => 12, 1 => 12514, 2 => 4695, 3 => 37190, 4 => 21379, 5 => 18723, 6 => 5802, 7 => 7182, 8 => 2529, 9 => 29936, 10 => 35860, 11 => 28338, 12 => 10835),
    14 => integer_vector_t'(0 => 12, 1 => 34283, 2 => 25610, 3 => 33026, 4 => 31017, 5 => 21259, 6 => 2165, 7 => 21807, 8 => 37578, 9 => 1175, 10 => 16710, 11 => 21939, 12 => 30841),
    15 => integer_vector_t'(0 => 12, 1 => 27292, 2 => 33730, 3 => 6836, 4 => 26476, 5 => 27539, 6 => 35784, 7 => 18245, 8 => 16394, 9 => 17939, 10 => 23094, 11 => 19216, 12 => 17432),
    16 => integer_vector_t'(0 => 12, 1 => 11655, 2 => 6183, 3 => 38708, 4 => 28408, 5 => 35157, 6 => 17089, 7 => 13998, 8 => 36029, 9 => 15052, 10 => 16617, 11 => 5638, 12 => 36464),
    17 => integer_vector_t'(0 => 12, 1 => 15693, 2 => 28923, 3 => 26245, 4 => 9432, 5 => 11675, 6 => 25720, 7 => 26405, 8 => 5838, 9 => 31851, 10 => 26898, 11 => 8090, 12 => 37037),
    18 => integer_vector_t'(0 => 12, 1 => 24418, 2 => 27583, 3 => 7959, 4 => 35562, 5 => 37771, 6 => 17784, 7 => 11382, 8 => 11156, 9 => 37855, 10 => 7073, 11 => 21685, 12 => 34515),
    19 => integer_vector_t'(0 => 12, 1 => 10977, 2 => 13633, 3 => 30969, 4 => 7516, 5 => 11943, 6 => 18199, 7 => 5231, 8 => 13825, 9 => 19589, 10 => 23661, 11 => 11150, 12 => 35602),
    20 => integer_vector_t'(0 => 12, 1 => 19124, 2 => 30774, 3 => 6670, 4 => 37344, 5 => 16510, 6 => 26317, 7 => 23518, 8 => 22957, 9 => 6348, 10 => 34069, 11 => 8845, 12 => 20175),
    21 => integer_vector_t'(0 => 12, 1 => 34985, 2 => 14441, 3 => 25668, 4 => 4116, 5 => 3019, 6 => 21049, 7 => 37308, 8 => 24551, 9 => 24727, 10 => 20104, 11 => 24850, 12 => 12114),
    22 => integer_vector_t'(0 => 12, 1 => 38187, 2 => 28527, 3 => 13108, 4 => 13985, 5 => 1425, 6 => 21477, 7 => 30807, 8 => 8613, 9 => 26241, 10 => 33368, 11 => 35913, 12 => 32477),
    23 => integer_vector_t'(0 => 12, 1 => 5903, 2 => 34390, 3 => 24641, 4 => 26556, 5 => 23007, 6 => 27305, 7 => 38247, 8 => 2621, 9 => 9122, 10 => 32806, 11 => 21554, 12 => 18685),
    24 => integer_vector_t'(0 => 3, 1 => 17287, 2 => 27292, 3 => 19033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25796, 2 => 31795, 3 => 12152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 12184, 2 => 35088, 3 => 31226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 38263, 2 => 33386, 3 => 24892, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 23114, 2 => 37995, 3 => 29796, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 34336, 2 => 10551, 3 => 36245, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 35407, 2 => 175, 3 => 7203, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 14654, 2 => 38201, 3 => 22605, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 28404, 2 => 6595, 3 => 1018, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 19932, 2 => 3524, 3 => 29305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 31749, 2 => 20247, 3 => 8128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 18026, 2 => 36357, 3 => 26735, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7543, 2 => 29767, 3 => 13588, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 13333, 2 => 25965, 3 => 8463, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 14504, 2 => 36796, 3 => 19710, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4528, 2 => 25299, 3 => 7318, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 35091, 2 => 25550, 3 => 14798, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 7824, 2 => 215, 3 => 1248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 30848, 2 => 5362, 3 => 17291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 28932, 2 => 30249, 3 => 27073, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 13062, 2 => 2103, 3 => 16206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 7129, 2 => 32062, 3 => 19612, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 9512, 2 => 21936, 3 => 38833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 35849, 2 => 33754, 3 => 23450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18705, 2 => 28656, 3 => 18111, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 22749, 2 => 27456, 3 => 32187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 28229, 2 => 31684, 3 => 30160, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15293, 2 => 8483, 3 => 28002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 14880, 2 => 13334, 3 => 12584, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 28646, 2 => 2558, 3 => 19687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 6259, 2 => 4499, 3 => 26336, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 11952, 2 => 28386, 3 => 8405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 10609, 2 => 961, 3 => 7582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 10423, 2 => 13191, 3 => 26818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 15922, 2 => 36654, 3 => 21450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 10492, 2 => 1532, 3 => 1205, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 30551, 2 => 36482, 3 => 22153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 5156, 2 => 11330, 3 => 34243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 28616, 2 => 35369, 3 => 13322, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 8962, 2 => 1485, 3 => 21186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 23541, 2 => 17445, 3 => 35561, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 33133, 2 => 11593, 3 => 19895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 33917, 2 => 7863, 3 => 33651, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 20063, 2 => 28331, 3 => 10702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 13195, 2 => 21107, 3 => 21859, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 4364, 2 => 31137, 3 => 4804, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 5585, 2 => 2037, 3 => 4830, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 30672, 2 => 16927, 3 => 14800, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_4.csv, table is 135x164 (2767.5 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_4 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 134)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 0, 2 => 6385, 3 => 7901, 4 => 14611, 5 => 13389, 6 => 11200, 7 => 3252, 8 => 5243, 9 => 2504, 10 => 2722, 11 => 821, 12 => 7374),
    1 => integer_vector_t'(0 => 12, 1 => 1, 2 => 11359, 3 => 2698, 4 => 357, 5 => 13824, 6 => 12772, 7 => 7244, 8 => 6752, 9 => 15310, 10 => 852, 11 => 2001, 12 => 11417),
    2 => integer_vector_t'(0 => 12, 1 => 2, 2 => 7862, 3 => 7977, 4 => 6321, 5 => 13612, 6 => 12197, 7 => 14449, 8 => 15137, 9 => 13860, 10 => 1708, 11 => 6399, 12 => 13444),
    3 => integer_vector_t'(0 => 12, 1 => 3, 2 => 1560, 3 => 11804, 4 => 6975, 5 => 13292, 6 => 3646, 7 => 3812, 8 => 8772, 9 => 7306, 10 => 5795, 11 => 14327, 12 => 7866),
    4 => integer_vector_t'(0 => 12, 1 => 4, 2 => 7626, 3 => 11407, 4 => 14599, 5 => 9689, 6 => 1628, 7 => 2113, 8 => 10809, 9 => 9283, 10 => 1230, 11 => 15241, 12 => 4870),
    5 => integer_vector_t'(0 => 12, 1 => 5, 2 => 1610, 3 => 5699, 4 => 15876, 5 => 9446, 6 => 12515, 7 => 1400, 8 => 6303, 9 => 5411, 10 => 14181, 11 => 13925, 12 => 7358),
    6 => integer_vector_t'(0 => 12, 1 => 6, 2 => 4059, 3 => 8836, 4 => 3405, 5 => 7853, 6 => 7992, 7 => 15336, 8 => 5970, 9 => 10368, 10 => 10278, 11 => 9675, 12 => 4651),
    7 => integer_vector_t'(0 => 12, 1 => 7, 2 => 4441, 3 => 3963, 4 => 9153, 5 => 2109, 6 => 12683, 7 => 7459, 8 => 12030, 9 => 12221, 10 => 629, 11 => 15212, 12 => 406),
    8 => integer_vector_t'(0 => 12, 1 => 8, 2 => 6007, 3 => 8411, 4 => 5771, 5 => 3497, 6 => 543, 7 => 14202, 8 => 875, 9 => 9186, 10 => 6235, 11 => 13908, 12 => 3563),
    9 => integer_vector_t'(0 => 12, 1 => 9, 2 => 3232, 3 => 6625, 4 => 4795, 5 => 546, 6 => 9781, 7 => 2071, 8 => 7312, 9 => 3399, 10 => 7250, 11 => 4932, 12 => 12652),
    10 => integer_vector_t'(0 => 12, 1 => 10, 2 => 8820, 3 => 10088, 4 => 11090, 5 => 7069, 6 => 6585, 7 => 13134, 8 => 10158, 9 => 7183, 10 => 488, 11 => 7455, 12 => 9238),
    11 => integer_vector_t'(0 => 12, 1 => 11, 2 => 1903, 3 => 10818, 4 => 119, 5 => 215, 6 => 7558, 7 => 11046, 8 => 10615, 9 => 11545, 10 => 14784, 11 => 7961, 12 => 15619),
    12 => integer_vector_t'(0 => 12, 1 => 12, 2 => 3655, 3 => 8736, 4 => 4917, 5 => 15874, 6 => 5129, 7 => 2134, 8 => 15944, 9 => 14768, 10 => 7150, 11 => 2692, 12 => 1469),
    13 => integer_vector_t'(0 => 12, 1 => 13, 2 => 8316, 3 => 3820, 4 => 505, 5 => 8923, 6 => 6757, 7 => 806, 8 => 7957, 9 => 4216, 10 => 15589, 11 => 13244, 12 => 2622),
    14 => integer_vector_t'(0 => 12, 1 => 14, 2 => 14463, 3 => 4852, 4 => 15733, 5 => 3041, 6 => 11193, 7 => 12860, 8 => 13673, 9 => 8152, 10 => 6551, 11 => 15108, 12 => 8758),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3149, 3 => 11981, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 13416, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 13098, 3 => 13352, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 2009, 3 => 14460, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 7207, 3 => 4314, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 3312, 3 => 3945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4418, 3 => 6248, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 2669, 3 => 13975, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 7571, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14172, 3 => 2967, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7271, 3 => 7138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6135, 3 => 13670, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 7490, 3 => 14559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8657, 3 => 2466, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8599, 3 => 12834, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 3470, 3 => 3152, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13917, 3 => 4365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 6024, 3 => 13730, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 10973, 3 => 14182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 2464, 3 => 13167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 5281, 3 => 15049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 36, 2 => 1103, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 37, 2 => 2058, 3 => 1069, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 38, 2 => 9654, 3 => 6095, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 39, 2 => 14311, 3 => 7667, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 40, 2 => 15617, 3 => 8146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 41, 2 => 4588, 3 => 11218, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 42, 2 => 13660, 3 => 6243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 43, 2 => 8578, 3 => 7874, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 44, 2 => 11741, 3 => 2686, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1022, 3 => 1264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 1, 2 => 12604, 3 => 9965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 2, 2 => 8217, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3156, 3 => 11793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 4, 2 => 354, 3 => 1514, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6978, 3 => 14058, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 6, 2 => 7922, 3 => 16079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 7, 2 => 15087, 3 => 12138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5053, 3 => 6470, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 9, 2 => 12687, 3 => 14932, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15458, 3 => 1763, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8121, 3 => 1721, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 12, 2 => 12431, 3 => 549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4129, 3 => 7091, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1426, 3 => 8415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9783, 3 => 7604, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6295, 3 => 11329, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1409, 3 => 12061, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 18, 2 => 8065, 3 => 9087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2918, 3 => 8438, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1293, 3 => 14115, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 21, 2 => 3922, 3 => 13851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3851, 3 => 4000, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5865, 3 => 1768, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2655, 3 => 14957, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 25, 2 => 5565, 3 => 6332, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4303, 3 => 12631, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11653, 3 => 12236, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 28, 2 => 16025, 3 => 7632, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4655, 3 => 14128, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 30, 2 => 9584, 3 => 13123, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 31, 2 => 13987, 3 => 9597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 32, 2 => 15409, 3 => 12110, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 33, 2 => 8754, 3 => 15490, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 34, 2 => 7416, 3 => 15325, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2909, 3 => 15549, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 36, 2 => 2995, 3 => 8257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 37, 2 => 9406, 3 => 4791, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 38, 2 => 11111, 3 => 4854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 39, 2 => 2812, 3 => 8521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 40, 2 => 8476, 3 => 14717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7820, 3 => 15360, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 42, 2 => 1179, 3 => 7939, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 43, 2 => 2357, 3 => 8678, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 44, 2 => 7703, 3 => 6216, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3477, 3 => 7067, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3931, 3 => 13845, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7675, 3 => 12899, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1754, 3 => 8187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7785, 3 => 1400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 9213, 3 => 5891, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2494, 3 => 7703, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2576, 3 => 7902, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4821, 3 => 15682, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 10426, 3 => 11935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1810, 3 => 904, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 11332, 3 => 9264, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11312, 3 => 3570, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 14916, 3 => 2650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7679, 3 => 7842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6089, 3 => 13084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3938, 3 => 2751, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8509, 3 => 4648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 12204, 3 => 8917, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5749, 3 => 12443, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12613, 3 => 4431, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1344, 3 => 4014, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 8488, 3 => 13850, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1730, 3 => 14896, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 14942, 3 => 7126, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 14983, 3 => 8863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6578, 3 => 8564, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 4947, 3 => 396, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 297, 3 => 12805, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 13878, 3 => 6692, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11857, 3 => 11186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 31, 2 => 14395, 3 => 11493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 32, 2 => 16145, 3 => 12251, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 33, 2 => 13462, 3 => 7428, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 34, 2 => 14526, 3 => 13119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 35, 2 => 2535, 3 => 11243, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 36, 2 => 6465, 3 => 12690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 37, 2 => 6872, 3 => 9334, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 38, 2 => 15371, 3 => 14023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 39, 2 => 8101, 3 => 10187, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 40, 2 => 11963, 3 => 4848, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 41, 2 => 15125, 3 => 6119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 42, 2 => 8051, 3 => 14465, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 43, 2 => 11139, 3 => 5167, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 44, 2 => 2883, 3 => 14521, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C3_5.csv, table is 108x184 (2484.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 15, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15, 9 => 15, 10 => 15, 11 => 15, 12 => 15);

  constant LDPC_TABLE_FECFRAME_NORMAL_C3_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 107)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 22422, 2 => 10282, 3 => 11626, 4 => 19997, 5 => 11161, 6 => 2922, 7 => 3122, 8 => 99, 9 => 5625, 10 => 17064, 11 => 8270, 12 => 179),
    1 => integer_vector_t'(0 => 12, 1 => 25087, 2 => 16218, 3 => 17015, 4 => 828, 5 => 20041, 6 => 25656, 7 => 4186, 8 => 11629, 9 => 22599, 10 => 17305, 11 => 22515, 12 => 6463),
    2 => integer_vector_t'(0 => 12, 1 => 11049, 2 => 22853, 3 => 25706, 4 => 14388, 5 => 5500, 6 => 19245, 7 => 8732, 8 => 2177, 9 => 13555, 10 => 11346, 11 => 17265, 12 => 3069),
    3 => integer_vector_t'(0 => 12, 1 => 16581, 2 => 22225, 3 => 12563, 4 => 19717, 5 => 23577, 6 => 11555, 7 => 25496, 8 => 6853, 9 => 25403, 10 => 5218, 11 => 15925, 12 => 21766),
    4 => integer_vector_t'(0 => 12, 1 => 16529, 2 => 14487, 3 => 7643, 4 => 10715, 5 => 17442, 6 => 11119, 7 => 5679, 8 => 14155, 9 => 24213, 10 => 21000, 11 => 1116, 12 => 15620),
    5 => integer_vector_t'(0 => 12, 1 => 5340, 2 => 8636, 3 => 16693, 4 => 1434, 5 => 5635, 6 => 6516, 7 => 9482, 8 => 20189, 9 => 1066, 10 => 15013, 11 => 25361, 12 => 14243),
    6 => integer_vector_t'(0 => 12, 1 => 18506, 2 => 22236, 3 => 20912, 4 => 8952, 5 => 5421, 6 => 15691, 7 => 6126, 8 => 21595, 9 => 500, 10 => 6904, 11 => 13059, 12 => 6802),
    7 => integer_vector_t'(0 => 12, 1 => 8433, 2 => 4694, 3 => 5524, 4 => 14216, 5 => 3685, 6 => 19721, 7 => 25420, 8 => 9937, 9 => 23813, 10 => 9047, 11 => 25651, 12 => 16826),
    8 => integer_vector_t'(0 => 12, 1 => 21500, 2 => 24814, 3 => 6344, 4 => 17382, 5 => 7064, 6 => 13929, 7 => 4004, 8 => 16552, 9 => 12818, 10 => 8720, 11 => 5286, 12 => 2206),
    9 => integer_vector_t'(0 => 12, 1 => 22517, 2 => 2429, 3 => 19065, 4 => 2921, 5 => 21611, 6 => 1873, 7 => 7507, 8 => 5661, 9 => 23006, 10 => 23128, 11 => 20543, 12 => 19777),
    10 => integer_vector_t'(0 => 12, 1 => 1770, 2 => 4636, 3 => 20900, 4 => 14931, 5 => 9247, 6 => 12340, 7 => 11008, 8 => 12966, 9 => 4471, 10 => 2731, 11 => 16445, 12 => 791),
    11 => integer_vector_t'(0 => 12, 1 => 6635, 2 => 14556, 3 => 18865, 4 => 22421, 5 => 22124, 6 => 12697, 7 => 9803, 8 => 25485, 9 => 7744, 10 => 18254, 11 => 11313, 12 => 9004),
    12 => integer_vector_t'(0 => 12, 1 => 19982, 2 => 23963, 3 => 18912, 4 => 7206, 5 => 12500, 6 => 4382, 7 => 20067, 8 => 6177, 9 => 21007, 10 => 1195, 11 => 23547, 12 => 24837),
    13 => integer_vector_t'(0 => 12, 1 => 756, 2 => 11158, 3 => 14646, 4 => 20534, 5 => 3647, 6 => 17728, 7 => 11676, 8 => 11843, 9 => 12937, 10 => 4402, 11 => 8261, 12 => 22944),
    14 => integer_vector_t'(0 => 12, 1 => 9306, 2 => 24009, 3 => 10012, 4 => 11081, 5 => 3746, 6 => 24325, 7 => 8060, 8 => 19826, 9 => 842, 10 => 8836, 11 => 2898, 12 => 5019),
    15 => integer_vector_t'(0 => 12, 1 => 7575, 2 => 7455, 3 => 25244, 4 => 4736, 5 => 14400, 6 => 22981, 7 => 5543, 8 => 8006, 9 => 24203, 10 => 13053, 11 => 1120, 12 => 5128),
    16 => integer_vector_t'(0 => 12, 1 => 3482, 2 => 9270, 3 => 13059, 4 => 15825, 5 => 7453, 6 => 23747, 7 => 3656, 8 => 24585, 9 => 16542, 10 => 17507, 11 => 22462, 12 => 14670),
    17 => integer_vector_t'(0 => 12, 1 => 15627, 2 => 15290, 3 => 4198, 4 => 22748, 5 => 5842, 6 => 13395, 7 => 23918, 8 => 16985, 9 => 14929, 10 => 3726, 11 => 25350, 12 => 24157),
    18 => integer_vector_t'(0 => 12, 1 => 24896, 2 => 16365, 3 => 16423, 4 => 13461, 5 => 16615, 6 => 8107, 7 => 24741, 8 => 3604, 9 => 25904, 10 => 8716, 11 => 9604, 12 => 20365),
    19 => integer_vector_t'(0 => 12, 1 => 3729, 2 => 17245, 3 => 18448, 4 => 9862, 5 => 20831, 6 => 25326, 7 => 20517, 8 => 24618, 9 => 13282, 10 => 5099, 11 => 14183, 12 => 8804),
    20 => integer_vector_t'(0 => 12, 1 => 16455, 2 => 17646, 3 => 15376, 4 => 18194, 5 => 25528, 6 => 1777, 7 => 6066, 8 => 21855, 9 => 14372, 10 => 12517, 11 => 4488, 12 => 17490),
    21 => integer_vector_t'(0 => 12, 1 => 1400, 2 => 8135, 3 => 23375, 4 => 20879, 5 => 8476, 6 => 4084, 7 => 12936, 8 => 25536, 9 => 22309, 10 => 16582, 11 => 6402, 12 => 24360),
    22 => integer_vector_t'(0 => 12, 1 => 25119, 2 => 23586, 3 => 128, 4 => 4761, 5 => 10443, 6 => 22536, 7 => 8607, 8 => 9752, 9 => 25446, 10 => 15053, 11 => 1856, 12 => 4040),
    23 => integer_vector_t'(0 => 12, 1 => 377, 2 => 21160, 3 => 13474, 4 => 5451, 5 => 17170, 6 => 5938, 7 => 10256, 8 => 11972, 9 => 24210, 10 => 17833, 11 => 22047, 12 => 16108),
    24 => integer_vector_t'(0 => 12, 1 => 13075, 2 => 9648, 3 => 24546, 4 => 13150, 5 => 23867, 6 => 7309, 7 => 19798, 8 => 2988, 9 => 16858, 10 => 4825, 11 => 23950, 12 => 15125),
    25 => integer_vector_t'(0 => 12, 1 => 20526, 2 => 3553, 3 => 11525, 4 => 23366, 5 => 2452, 6 => 17626, 7 => 19265, 8 => 20172, 9 => 18060, 10 => 24593, 11 => 13255, 12 => 1552),
    26 => integer_vector_t'(0 => 12, 1 => 18839, 2 => 21132, 3 => 20119, 4 => 15214, 5 => 14705, 6 => 7096, 7 => 10174, 8 => 5663, 9 => 18651, 10 => 19700, 11 => 12524, 12 => 14033),
    27 => integer_vector_t'(0 => 12, 1 => 4127, 2 => 2971, 3 => 17499, 4 => 16287, 5 => 22368, 6 => 21463, 7 => 7943, 8 => 18880, 9 => 5567, 10 => 8047, 11 => 23363, 12 => 6797),
    28 => integer_vector_t'(0 => 12, 1 => 10651, 2 => 24471, 3 => 14325, 4 => 4081, 5 => 7258, 6 => 4949, 7 => 7044, 8 => 1078, 9 => 797, 10 => 22910, 11 => 20474, 12 => 4318),
    29 => integer_vector_t'(0 => 12, 1 => 21374, 2 => 13231, 3 => 22985, 4 => 5056, 5 => 3821, 6 => 23718, 7 => 14178, 8 => 9978, 9 => 19030, 10 => 23594, 11 => 8895, 12 => 25358),
    30 => integer_vector_t'(0 => 12, 1 => 6199, 2 => 22056, 3 => 7749, 4 => 13310, 5 => 3999, 6 => 23697, 7 => 16445, 8 => 22636, 9 => 5225, 10 => 22437, 11 => 24153, 12 => 9442),
    31 => integer_vector_t'(0 => 12, 1 => 7978, 2 => 12177, 3 => 2893, 4 => 20778, 5 => 3175, 6 => 8645, 7 => 11863, 8 => 24623, 9 => 10311, 10 => 25767, 11 => 17057, 12 => 3691),
    32 => integer_vector_t'(0 => 12, 1 => 20473, 2 => 11294, 3 => 9914, 4 => 22815, 5 => 2574, 6 => 8439, 7 => 3699, 8 => 5431, 9 => 24840, 10 => 21908, 11 => 16088, 12 => 18244),
    33 => integer_vector_t'(0 => 12, 1 => 8208, 2 => 5755, 3 => 19059, 4 => 8541, 5 => 24924, 6 => 6454, 7 => 11234, 8 => 10492, 9 => 16406, 10 => 10831, 11 => 11436, 12 => 9649),
    34 => integer_vector_t'(0 => 12, 1 => 16264, 2 => 11275, 3 => 24953, 4 => 2347, 5 => 12667, 6 => 19190, 7 => 7257, 8 => 7174, 9 => 24819, 10 => 2938, 11 => 2522, 12 => 11749),
    35 => integer_vector_t'(0 => 12, 1 => 3627, 2 => 5969, 3 => 13862, 4 => 1538, 5 => 23176, 6 => 6353, 7 => 2855, 8 => 17720, 9 => 2472, 10 => 7428, 11 => 573, 12 => 15036),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 18539, 3 => 18661, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 10502, 3 => 3002, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 9368, 3 => 10761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 12299, 3 => 7828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 15048, 3 => 13362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 18444, 3 => 24640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 20775, 3 => 19175, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 18970, 3 => 10971, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5329, 3 => 19982, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 11296, 3 => 18655, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 15046, 3 => 20659, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 7300, 3 => 22140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 22029, 3 => 14477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 11129, 3 => 742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 13254, 3 => 13813, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 19234, 3 => 13273, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6079, 3 => 21122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 22782, 3 => 5828, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 19775, 3 => 4247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1660, 3 => 19413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4403, 3 => 3649, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 13371, 3 => 25851, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 22770, 3 => 21784, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 10757, 3 => 14131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 16071, 3 => 21617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 6393, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 597, 3 => 19968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5743, 3 => 8084, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 6770, 3 => 9548, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 4285, 3 => 17542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 13568, 3 => 22599, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 1786, 3 => 4617, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 23238, 3 => 11648, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 19627, 3 => 2030, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 13601, 3 => 13458, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 13740, 3 => 17328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 36, 2 => 25012, 3 => 13944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 37, 2 => 22513, 3 => 6687, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 38, 2 => 4934, 3 => 12587, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 39, 2 => 21197, 3 => 5133, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 40, 2 => 22705, 3 => 6938, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 41, 2 => 7534, 3 => 24633, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 42, 2 => 24400, 3 => 12797, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 43, 2 => 21911, 3 => 25712, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 44, 2 => 12039, 3 => 1140, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 45, 2 => 24306, 3 => 1021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 46, 2 => 14012, 3 => 20747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 47, 2 => 11265, 3 => 15219, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 48, 2 => 4670, 3 => 15531, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 49, 2 => 9417, 3 => 14359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 50, 2 => 2415, 3 => 6504, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 51, 2 => 24964, 3 => 24690, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 52, 2 => 14443, 3 => 8816, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 53, 2 => 6926, 3 => 1291, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 54, 2 => 6209, 3 => 20806, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 55, 2 => 13915, 3 => 4079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 56, 2 => 24410, 3 => 13196, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 57, 2 => 13505, 3 => 6117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 58, 2 => 9869, 3 => 8220, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 59, 2 => 1570, 3 => 6044, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 60, 2 => 25780, 3 => 17387, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 61, 2 => 20671, 3 => 24913, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 62, 2 => 24558, 3 => 20591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 63, 2 => 12402, 3 => 3702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 64, 2 => 8314, 3 => 1357, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 65, 2 => 20071, 3 => 14616, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 66, 2 => 17014, 3 => 3688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 67, 2 => 19837, 3 => 946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 68, 2 => 15195, 3 => 12136, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 69, 2 => 7758, 3 => 22808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 70, 2 => 3564, 3 => 2925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 71, 2 => 3434, 3 => 7769, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C4_5.csv, table is 144x150 (2700.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C4_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 143)(0 to 11)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 11, 1 => 0, 2 => 149, 3 => 11212, 4 => 5575, 5 => 6360, 6 => 12559, 7 => 8108, 8 => 8505, 9 => 408, 10 => 10026, 11 => 12828),
    1 => integer_vector_t'(0 => 11, 1 => 1, 2 => 5237, 3 => 490, 4 => 10677, 5 => 4998, 6 => 3869, 7 => 3734, 8 => 3092, 9 => 3509, 10 => 7703, 11 => 10305),
    2 => integer_vector_t'(0 => 11, 1 => 2, 2 => 8742, 3 => 5553, 4 => 2820, 5 => 7085, 6 => 12116, 7 => 10485, 8 => 564, 9 => 7795, 10 => 2972, 11 => 2157),
    3 => integer_vector_t'(0 => 11, 1 => 3, 2 => 2699, 3 => 4304, 4 => 8350, 5 => 712, 6 => 2841, 7 => 3250, 8 => 4731, 9 => 10105, 10 => 517, 11 => 7516),
    4 => integer_vector_t'(0 => 11, 1 => 4, 2 => 12067, 3 => 1351, 4 => 11992, 5 => 12191, 6 => 11267, 7 => 5161, 8 => 537, 9 => 6166, 10 => 4246, 11 => 2363),
    5 => integer_vector_t'(0 => 11, 1 => 5, 2 => 6828, 3 => 7107, 4 => 2127, 5 => 3724, 6 => 5743, 7 => 11040, 8 => 10756, 9 => 4073, 10 => 1011, 11 => 3422),
    6 => integer_vector_t'(0 => 11, 1 => 6, 2 => 11259, 3 => 1216, 4 => 9526, 5 => 1466, 6 => 10816, 7 => 940, 8 => 3744, 9 => 2815, 10 => 11506, 11 => 11573),
    7 => integer_vector_t'(0 => 11, 1 => 7, 2 => 4549, 3 => 11507, 4 => 1118, 5 => 1274, 6 => 11751, 7 => 5207, 8 => 7854, 9 => 12803, 10 => 4047, 11 => 6484),
    8 => integer_vector_t'(0 => 11, 1 => 8, 2 => 8430, 3 => 4115, 4 => 9440, 5 => 413, 6 => 4455, 7 => 2262, 8 => 7915, 9 => 12402, 10 => 8579, 11 => 7052),
    9 => integer_vector_t'(0 => 11, 1 => 9, 2 => 3885, 3 => 9126, 4 => 5665, 5 => 4505, 6 => 2343, 7 => 253, 8 => 4707, 9 => 3742, 10 => 4166, 11 => 1556),
    10 => integer_vector_t'(0 => 11, 1 => 10, 2 => 1704, 3 => 8936, 4 => 6775, 5 => 8639, 6 => 8179, 7 => 7954, 8 => 8234, 9 => 7850, 10 => 8883, 11 => 8713),
    11 => integer_vector_t'(0 => 11, 1 => 11, 2 => 11716, 3 => 4344, 4 => 9087, 5 => 11264, 6 => 2274, 7 => 8832, 8 => 9147, 9 => 11930, 10 => 6054, 11 => 5455),
    12 => integer_vector_t'(0 => 11, 1 => 12, 2 => 7323, 3 => 3970, 4 => 10329, 5 => 2170, 6 => 8262, 7 => 3854, 8 => 2087, 9 => 12899, 10 => 9497, 11 => 11700),
    13 => integer_vector_t'(0 => 11, 1 => 13, 2 => 4418, 3 => 1467, 4 => 2490, 5 => 5841, 6 => 817, 7 => 11453, 8 => 533, 9 => 11217, 10 => 11962, 11 => 5251),
    14 => integer_vector_t'(0 => 11, 1 => 14, 2 => 1541, 3 => 4525, 4 => 7976, 5 => 3457, 6 => 9536, 7 => 7725, 8 => 3788, 9 => 2982, 10 => 6307, 11 => 5997),
    15 => integer_vector_t'(0 => 11, 1 => 15, 2 => 11484, 3 => 2739, 4 => 4023, 5 => 12107, 6 => 6516, 7 => 551, 8 => 2572, 9 => 6628, 10 => 8150, 11 => 9852),
    16 => integer_vector_t'(0 => 11, 1 => 16, 2 => 6070, 3 => 1761, 4 => 4627, 5 => 6534, 6 => 7913, 7 => 3730, 8 => 11866, 9 => 1813, 10 => 12306, 11 => 8249),
    17 => integer_vector_t'(0 => 11, 1 => 17, 2 => 12441, 3 => 5489, 4 => 8748, 5 => 7837, 6 => 7660, 7 => 2102, 8 => 11341, 9 => 2936, 10 => 6712, 11 => 11977),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10155, 3 => 4210, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1010, 3 => 10483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 8900, 3 => 10250, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 10243, 3 => 12278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 7070, 3 => 4397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 12271, 3 => 3887, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 11980, 3 => 6836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 9514, 3 => 4356, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 7137, 3 => 10281, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 11881, 3 => 2526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 1969, 3 => 11477, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3044, 3 => 10921, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 30, 2 => 2236, 3 => 8724, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9104, 3 => 6340, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 32, 2 => 7342, 3 => 8582, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 33, 2 => 11675, 3 => 10405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 34, 2 => 6467, 3 => 12775, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 35, 2 => 3186, 3 => 12198, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 9621, 3 => 11445, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7486, 3 => 5611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4319, 3 => 4879, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2196, 3 => 344, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 7527, 3 => 6650, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 10693, 3 => 2440, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6755, 3 => 2706, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5144, 3 => 5998, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 11043, 3 => 8033, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4846, 3 => 4435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4157, 3 => 9228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 12270, 3 => 6562, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 11954, 3 => 7592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 7420, 3 => 2592, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 8810, 3 => 9636, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 689, 3 => 5430, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 920, 3 => 1304, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1253, 3 => 11934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9559, 3 => 6016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 19, 2 => 312, 3 => 7589, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4439, 3 => 4197, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4002, 3 => 9555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12232, 3 => 7779, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 23, 2 => 1494, 3 => 8782, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 24, 2 => 10749, 3 => 3969, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4368, 3 => 3479, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6316, 3 => 5342, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2455, 3 => 3493, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12157, 3 => 7405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 29, 2 => 6598, 3 => 11495, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 30, 2 => 11805, 3 => 4455, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9625, 3 => 2090, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 32, 2 => 4731, 3 => 2321, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 33, 2 => 3578, 3 => 2608, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 34, 2 => 8504, 3 => 1849, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 35, 2 => 4027, 3 => 1151, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5647, 3 => 4935, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4219, 3 => 1870, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10968, 3 => 8054, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6970, 3 => 5447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3217, 3 => 5638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 8972, 3 => 669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5618, 3 => 12472, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1457, 3 => 1280, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 8868, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8866, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 8371, 3 => 5972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 266, 3 => 4405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3706, 3 => 3244, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 6039, 3 => 5844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7200, 3 => 3283, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1502, 3 => 11282, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 12318, 3 => 2202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4523, 3 => 965, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 18, 2 => 9587, 3 => 7011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 19, 2 => 2552, 3 => 2051, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 20, 2 => 12045, 3 => 10306, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 21, 2 => 11070, 3 => 5104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6627, 3 => 6906, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 23, 2 => 9889, 3 => 2121, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 24, 2 => 829, 3 => 9701, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2201, 3 => 1819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6689, 3 => 12925, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 27, 2 => 2139, 3 => 8757, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12004, 3 => 5948, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8704, 3 => 3191, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 30, 2 => 8171, 3 => 10933, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 31, 2 => 6297, 3 => 7116, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 32, 2 => 616, 3 => 7146, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 33, 2 => 5142, 3 => 9761, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 34, 2 => 10377, 3 => 8138, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7616, 3 => 5811, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7285, 3 => 9863, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 7764, 3 => 10867, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 12343, 3 => 9019, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4414, 3 => 8331, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3464, 3 => 642, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6960, 3 => 2039, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 786, 3 => 3021, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 710, 3 => 2086, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 7423, 3 => 5601, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 8120, 3 => 4885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 12385, 3 => 11990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9739, 3 => 10034, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 424, 3 => 10162, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1347, 3 => 7597, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1450, 3 => 112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 7965, 3 => 8478, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8945, 3 => 7397, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 6590, 3 => 8316, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6838, 3 => 9011, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6174, 3 => 9410, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 20, 2 => 255, 3 => 113, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 21, 2 => 6197, 3 => 5835, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 22, 2 => 12902, 3 => 3844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 23, 2 => 4377, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 24, 2 => 5478, 3 => 8672, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 25, 2 => 4453, 3 => 2132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 26, 2 => 9724, 3 => 1380, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 27, 2 => 12131, 3 => 11526, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 28, 2 => 12323, 3 => 9511, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 29, 2 => 8231, 3 => 1752, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 30, 2 => 497, 3 => 9022, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 31, 2 => 9288, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 32, 2 => 2481, 3 => 7515, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 33, 2 => 2696, 3 => 268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 34, 2 => 4023, 3 => 12341, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 35, 2 => 7108, 3 => 5553, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C5_6.csv, table is 150x177 (3318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 5, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14, 13 => 14);

  constant LDPC_TABLE_FECFRAME_NORMAL_C5_6 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 149)(0 to 13)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 4362, 3 => 416, 4 => 8909, 5 => 4156, 6 => 3216, 7 => 3112, 8 => 2560, 9 => 2912, 10 => 6405, 11 => 8593, 12 => 4969, 13 => 6723),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 2479, 3 => 1786, 4 => 8978, 5 => 3011, 6 => 4339, 7 => 9313, 8 => 6397, 9 => 2957, 10 => 7288, 11 => 5484, 12 => 6031, 13 => 10217),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 10175, 3 => 9009, 4 => 9889, 5 => 3091, 6 => 4985, 7 => 7267, 8 => 4092, 9 => 8874, 10 => 5671, 11 => 2777, 12 => 2189, 13 => 8716),
    3 => integer_vector_t'(0 => 13, 1 => 3, 2 => 9052, 3 => 4795, 4 => 3924, 5 => 3370, 6 => 10058, 7 => 1128, 8 => 9996, 9 => 10165, 10 => 9360, 11 => 4297, 12 => 434, 13 => 5138),
    4 => integer_vector_t'(0 => 13, 1 => 4, 2 => 2379, 3 => 7834, 4 => 4835, 5 => 2327, 6 => 9843, 7 => 804, 8 => 329, 9 => 8353, 10 => 7167, 11 => 3070, 12 => 1528, 13 => 7311),
    5 => integer_vector_t'(0 => 13, 1 => 5, 2 => 3435, 3 => 7871, 4 => 348, 5 => 3693, 6 => 1876, 7 => 6585, 8 => 10340, 9 => 7144, 10 => 5870, 11 => 2084, 12 => 4052, 13 => 2780),
    6 => integer_vector_t'(0 => 13, 1 => 6, 2 => 3917, 3 => 3111, 4 => 3476, 5 => 1304, 6 => 10331, 7 => 5939, 8 => 5199, 9 => 1611, 10 => 1991, 11 => 699, 12 => 8316, 13 => 9960),
    7 => integer_vector_t'(0 => 13, 1 => 7, 2 => 6883, 3 => 3237, 4 => 1717, 5 => 10752, 6 => 7891, 7 => 9764, 8 => 4745, 9 => 3888, 10 => 10009, 11 => 4176, 12 => 4614, 13 => 1567),
    8 => integer_vector_t'(0 => 13, 1 => 8, 2 => 10587, 3 => 2195, 4 => 1689, 5 => 2968, 6 => 5420, 7 => 2580, 8 => 2883, 9 => 6496, 10 => 111, 11 => 6023, 12 => 1024, 13 => 4449),
    9 => integer_vector_t'(0 => 13, 1 => 9, 2 => 3786, 3 => 8593, 4 => 2074, 5 => 3321, 6 => 5057, 7 => 1450, 8 => 3840, 9 => 5444, 10 => 6572, 11 => 3094, 12 => 9892, 13 => 1512),
    10 => integer_vector_t'(0 => 13, 1 => 10, 2 => 8548, 3 => 1848, 4 => 10372, 5 => 4585, 6 => 7313, 7 => 6536, 8 => 6379, 9 => 1766, 10 => 9462, 11 => 2456, 12 => 5606, 13 => 9975),
    11 => integer_vector_t'(0 => 13, 1 => 11, 2 => 8204, 3 => 10593, 4 => 7935, 5 => 3636, 6 => 3882, 7 => 394, 8 => 5968, 9 => 8561, 10 => 2395, 11 => 7289, 12 => 9267, 13 => 9978),
    12 => integer_vector_t'(0 => 13, 1 => 12, 2 => 7795, 3 => 74, 4 => 1633, 5 => 9542, 6 => 6867, 7 => 7352, 8 => 6417, 9 => 7568, 10 => 10623, 11 => 725, 12 => 2531, 13 => 9115),
    13 => integer_vector_t'(0 => 13, 1 => 13, 2 => 7151, 3 => 2482, 4 => 4260, 5 => 5003, 6 => 10105, 7 => 7419, 8 => 9203, 9 => 6691, 10 => 8798, 11 => 2092, 12 => 8263, 13 => 3755),
    14 => integer_vector_t'(0 => 13, 1 => 14, 2 => 3600, 3 => 570, 4 => 4527, 5 => 200, 6 => 9718, 7 => 6771, 8 => 1995, 9 => 8902, 10 => 5446, 11 => 768, 12 => 1103, 13 => 6520),
    15 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6304, 3 => 7621, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6498, 3 => 9209, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 17, 2 => 7293, 3 => 6786, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5950, 3 => 1708, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8521, 3 => 1793, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 20, 2 => 6174, 3 => 7854, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9773, 3 => 1190, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9517, 3 => 10268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2181, 3 => 9349, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 24, 2 => 1949, 3 => 5560, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 25, 2 => 1556, 3 => 555, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8600, 3 => 3827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 27, 2 => 5072, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7928, 3 => 3542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 29, 2 => 3226, 3 => 3762, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 7045, 3 => 2420, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 9645, 3 => 2641, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2774, 3 => 2452, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5331, 3 => 2031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 9400, 3 => 7503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1850, 3 => 2338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10456, 3 => 9774, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1692, 3 => 9276, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 8, 2 => 10037, 3 => 4038, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3964, 3 => 338, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 10, 2 => 2640, 3 => 5087, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 11, 2 => 858, 3 => 3473, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5582, 3 => 5683, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9523, 3 => 916, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4107, 3 => 1559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4506, 3 => 3491, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 16, 2 => 8191, 3 => 4182, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 17, 2 => 10192, 3 => 6157, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5668, 3 => 3305, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3449, 3 => 1540, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4766, 3 => 2697, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 21, 2 => 4069, 3 => 6675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 22, 2 => 1117, 3 => 1016, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5619, 3 => 3085, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 24, 2 => 8483, 3 => 8400, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 25, 2 => 8255, 3 => 394, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 26, 2 => 6338, 3 => 5042, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 27, 2 => 6174, 3 => 5119, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 28, 2 => 7203, 3 => 1989, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 29, 2 => 1781, 3 => 5174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1464, 3 => 3559, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3376, 3 => 4214, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 7238, 3 => 67, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 10595, 3 => 8831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1221, 3 => 6513, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5300, 3 => 4652, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1429, 3 => 9749, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7878, 3 => 5131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4435, 3 => 10284, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6331, 3 => 5507, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6662, 3 => 4941, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 9614, 3 => 10238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 8400, 3 => 8025, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 9156, 3 => 5630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7067, 3 => 8878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 9027, 3 => 3415, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1690, 3 => 3866, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2854, 3 => 8469, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6206, 3 => 630, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 363, 3 => 5453, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 20, 2 => 4125, 3 => 7008, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 21, 2 => 1612, 3 => 6702, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 22, 2 => 9069, 3 => 9226, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 23, 2 => 5767, 3 => 4060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 24, 2 => 3743, 3 => 9237, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 25, 2 => 7018, 3 => 5572, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 26, 2 => 8892, 3 => 4536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 27, 2 => 853, 3 => 6064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 28, 2 => 8069, 3 => 5893, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 29, 2 => 2051, 3 => 2885, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 10691, 3 => 3153, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3602, 3 => 4055, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 328, 3 => 1717, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 2219, 3 => 9299, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1939, 3 => 7898, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 617, 3 => 206, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 8544, 3 => 1374, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 10676, 3 => 3240, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6672, 3 => 9489, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3170, 3 => 7457, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7868, 3 => 5731, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6121, 3 => 10732, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4843, 3 => 9132, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 580, 3 => 9591, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 6267, 3 => 9290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3009, 3 => 2268, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 195, 3 => 2419, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 8016, 3 => 1557, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1516, 3 => 9195, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8062, 3 => 9064, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 20, 2 => 2095, 3 => 8968, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 21, 2 => 753, 3 => 7326, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 22, 2 => 6291, 3 => 3833, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2614, 3 => 7844, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 24, 2 => 2303, 3 => 646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 25, 2 => 2075, 3 => 611, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4687, 3 => 362, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 27, 2 => 8684, 3 => 9940, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4830, 3 => 2065, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7038, 3 => 1363, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1769, 3 => 7837, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3801, 3 => 1689, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 10070, 3 => 2359, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3667, 3 => 9918, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1914, 3 => 6920, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4244, 3 => 5669, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 10245, 3 => 7821, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7648, 3 => 3944, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3310, 3 => 5488, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 6346, 3 => 9666, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 7088, 3 => 6122, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1291, 3 => 7827, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 10592, 3 => 8945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3609, 3 => 7120, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 9168, 3 => 9112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6203, 3 => 8052, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3330, 3 => 2895, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4264, 3 => 10563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 10556, 3 => 6496, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 8807, 3 => 7645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 20, 2 => 1999, 3 => 4530, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 21, 2 => 9202, 3 => 6818, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 22, 2 => 3403, 3 => 1734, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 23, 2 => 2106, 3 => 9023, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 24, 2 => 6881, 3 => 3883, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 25, 2 => 3895, 3 => 2171, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 26, 2 => 4062, 3 => 6424, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 27, 2 => 3755, 3 => 9536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 28, 2 => 4683, 3 => 2131, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 29, 2 => 7347, 3 => 8027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C8_9.csv, table is 160x46 (920.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C8_9 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 159)(0 to 4)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 6235, 3 => 2848, 4 => 3222),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5800, 3 => 3492, 4 => 5348),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2757, 3 => 927, 4 => 90),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6961, 3 => 4516, 4 => 4739),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1172, 3 => 3237, 4 => 6264),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1927, 3 => 2425, 4 => 3683),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3714, 3 => 6309, 4 => 2495),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 3070, 3 => 6342, 4 => 7154),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2428, 3 => 613, 4 => 3761),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 2906, 3 => 264, 4 => 5927),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 1716, 3 => 1950, 4 => 4273),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4613, 3 => 6179, 4 => 3491),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 4865, 3 => 3286, 4 => 6005),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1343, 3 => 5923, 4 => 3529),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 4589, 3 => 4035, 4 => 2132),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 1579, 3 => 3920, 4 => 6737),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1644, 3 => 1191, 4 => 5998),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 1482, 3 => 2381, 4 => 4620),
    18 => integer_vector_t'(0 => 4, 1 => 18, 2 => 6791, 3 => 6014, 4 => 6596),
    19 => integer_vector_t'(0 => 4, 1 => 19, 2 => 2738, 3 => 5918, 4 => 3786),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5156, 3 => 6166, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1504, 3 => 4356, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 130, 3 => 1904, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 6027, 3 => 3187, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6718, 3 => 759, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 5, 2 => 6240, 3 => 2870, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2343, 3 => 1311, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1039, 3 => 5465, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 8, 2 => 6617, 3 => 2513, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1588, 3 => 5222, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 10, 2 => 6561, 3 => 535, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4765, 3 => 2054, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 12, 2 => 5966, 3 => 6892, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1969, 3 => 3869, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3571, 3 => 2420, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4632, 3 => 981, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3215, 3 => 4163, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 17, 2 => 973, 3 => 3117, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 18, 2 => 3802, 3 => 6198, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 19, 2 => 3794, 3 => 3948, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3196, 3 => 6126, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 1, 2 => 573, 3 => 1909, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 2, 2 => 850, 3 => 4034, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5622, 3 => 1601, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6005, 3 => 524, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5251, 3 => 5783, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 6, 2 => 172, 3 => 2032, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1875, 3 => 2475, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 8, 2 => 497, 3 => 1291, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2566, 3 => 3430, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1249, 3 => 740, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2944, 3 => 1948, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6528, 3 => 2899, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2243, 3 => 3616, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 14, 2 => 867, 3 => 3733, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1374, 3 => 4702, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4698, 3 => 2285, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4760, 3 => 3917, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1859, 3 => 4058, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6141, 3 => 3527, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2148, 3 => 5066, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1306, 3 => 145, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2319, 3 => 871, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3463, 3 => 1061, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5554, 3 => 6647, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5837, 3 => 339, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5821, 3 => 4932, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6356, 3 => 4756, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3930, 3 => 418, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 9, 2 => 211, 3 => 3094, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1007, 3 => 4928, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3584, 3 => 1235, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6982, 3 => 2869, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1612, 3 => 1013, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 14, 2 => 953, 3 => 4964, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4555, 3 => 4410, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4925, 3 => 4842, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5778, 3 => 600, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 18, 2 => 6509, 3 => 2417, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1260, 3 => 4903, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3369, 3 => 3031, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3557, 3 => 3224, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3028, 3 => 583, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3258, 3 => 440, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 4, 2 => 6226, 3 => 6655, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4895, 3 => 1094, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1481, 3 => 6847, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4433, 3 => 1932, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2107, 3 => 1649, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2119, 3 => 2065, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4003, 3 => 6388, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6720, 3 => 3622, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3694, 3 => 4521, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1164, 3 => 7050, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1965, 3 => 3613, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4331, 3 => 66, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2970, 3 => 1796, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4652, 3 => 3218, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 18, 2 => 1762, 3 => 4777, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 19, 2 => 5736, 3 => 1399, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 0, 2 => 970, 3 => 2572, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2062, 3 => 6599, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4597, 3 => 4870, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1228, 3 => 6913, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4159, 3 => 1037, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2916, 3 => 2362, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 6, 2 => 395, 3 => 1226, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6911, 3 => 4548, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4618, 3 => 2241, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4120, 3 => 4280, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5825, 3 => 474, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2154, 3 => 5558, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3793, 3 => 5471, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5707, 3 => 1595, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1403, 3 => 325, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6601, 3 => 5183, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6369, 3 => 4569, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4846, 3 => 896, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 18, 2 => 7092, 3 => 6184, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6764, 3 => 7127, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6358, 3 => 1951, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3117, 3 => 6960, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2710, 3 => 7062, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1133, 3 => 3604, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3694, 3 => 657, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1355, 3 => 110, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3329, 3 => 6736, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2505, 3 => 3407, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2462, 3 => 4806, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4216, 3 => 214, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5348, 3 => 5619, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 11, 2 => 6627, 3 => 6243, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 12, 2 => 2644, 3 => 5073, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 13, 2 => 4212, 3 => 5088, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3463, 3 => 3889, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5306, 3 => 478, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 16, 2 => 4320, 3 => 6121, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3961, 3 => 1125, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5699, 3 => 1195, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 19, 2 => 6511, 3 => 792, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3934, 3 => 2778, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3238, 3 => 6587, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1111, 3 => 6596, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1457, 3 => 6226, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1446, 3 => 3885, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3907, 3 => 4043, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6839, 3 => 2873, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1733, 3 => 5615, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5202, 3 => 4269, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3024, 3 => 4722, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5445, 3 => 6372, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 11, 2 => 370, 3 => 1828, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 12, 2 => 4695, 3 => 1600, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 13, 2 => 680, 3 => 2074, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1801, 3 => 6690, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2669, 3 => 1377, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 16, 2 => 2463, 3 => 1681, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 17, 2 => 5972, 3 => 5171, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 18, 2 => 5728, 3 => 4284, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 19, 2 => 1696, 3 => 1459, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_NORMAL_C9_10.csv, table is 162x46 (931.5 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant LDPC_TABLE_FECFRAME_NORMAL_C9_10 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 161)(0 to 4)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 5611, 3 => 2563, 4 => 2900),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 5220, 3 => 3143, 4 => 4813),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 2481, 3 => 834, 4 => 81),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 6265, 3 => 4064, 4 => 4265),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 1055, 3 => 2914, 4 => 5638),
    5 => integer_vector_t'(0 => 4, 1 => 5, 2 => 1734, 3 => 2182, 4 => 3315),
    6 => integer_vector_t'(0 => 4, 1 => 6, 2 => 3342, 3 => 5678, 4 => 2246),
    7 => integer_vector_t'(0 => 4, 1 => 7, 2 => 2185, 3 => 552, 4 => 3385),
    8 => integer_vector_t'(0 => 4, 1 => 8, 2 => 2615, 3 => 236, 4 => 5334),
    9 => integer_vector_t'(0 => 4, 1 => 9, 2 => 1546, 3 => 1755, 4 => 3846),
    10 => integer_vector_t'(0 => 4, 1 => 10, 2 => 4154, 3 => 5561, 4 => 3142),
    11 => integer_vector_t'(0 => 4, 1 => 11, 2 => 4382, 3 => 2957, 4 => 5400),
    12 => integer_vector_t'(0 => 4, 1 => 12, 2 => 1209, 3 => 5329, 4 => 3179),
    13 => integer_vector_t'(0 => 4, 1 => 13, 2 => 1421, 3 => 3528, 4 => 6063),
    14 => integer_vector_t'(0 => 4, 1 => 14, 2 => 1480, 3 => 1072, 4 => 5398),
    15 => integer_vector_t'(0 => 4, 1 => 15, 2 => 3843, 3 => 1777, 4 => 4369),
    16 => integer_vector_t'(0 => 4, 1 => 16, 2 => 1334, 3 => 2145, 4 => 4163),
    17 => integer_vector_t'(0 => 4, 1 => 17, 2 => 2368, 3 => 5055, 4 => 260),
    18 => integer_vector_t'(0 => 3, 1 => 0, 2 => 6118, 3 => 5405, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2994, 3 => 4370, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 2, 2 => 3405, 3 => 1669, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4640, 3 => 5550, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1354, 3 => 3921, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 5, 2 => 117, 3 => 1713, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 6, 2 => 5425, 3 => 2866, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 7, 2 => 6047, 3 => 683, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5616, 3 => 2582, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2108, 3 => 1179, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 10, 2 => 933, 3 => 4921, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5953, 3 => 2261, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1430, 3 => 4699, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5905, 3 => 480, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 14, 2 => 4289, 3 => 1846, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5374, 3 => 6208, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1775, 3 => 3476, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3216, 3 => 2178, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4165, 3 => 884, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2896, 3 => 3744, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 2801, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3423, 3 => 5579, 4 => -1),
    40 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3404, 3 => 3552, 4 => -1),
    41 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2876, 3 => 5515, 4 => -1),
    42 => integer_vector_t'(0 => 3, 1 => 6, 2 => 516, 3 => 1719, 4 => -1),
    43 => integer_vector_t'(0 => 3, 1 => 7, 2 => 765, 3 => 3631, 4 => -1),
    44 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5059, 3 => 1441, 4 => -1),
    45 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5629, 3 => 598, 4 => -1),
    46 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5405, 3 => 473, 4 => -1),
    47 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4724, 3 => 5210, 4 => -1),
    48 => integer_vector_t'(0 => 3, 1 => 12, 2 => 155, 3 => 1832, 4 => -1),
    49 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1689, 3 => 2229, 4 => -1),
    50 => integer_vector_t'(0 => 3, 1 => 14, 2 => 449, 3 => 1164, 4 => -1),
    51 => integer_vector_t'(0 => 3, 1 => 15, 2 => 2308, 3 => 3088, 4 => -1),
    52 => integer_vector_t'(0 => 3, 1 => 16, 2 => 1122, 3 => 669, 4 => -1),
    53 => integer_vector_t'(0 => 3, 1 => 17, 2 => 2268, 3 => 5758, 4 => -1),
    54 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5878, 3 => 2609, 4 => -1),
    55 => integer_vector_t'(0 => 3, 1 => 1, 2 => 782, 3 => 3359, 4 => -1),
    56 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1231, 3 => 4231, 4 => -1),
    57 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4225, 3 => 2052, 4 => -1),
    58 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4286, 3 => 3517, 4 => -1),
    59 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5531, 3 => 3184, 4 => -1),
    60 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1935, 3 => 4560, 4 => -1),
    61 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1174, 3 => 131, 4 => -1),
    62 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3115, 3 => 956, 4 => -1),
    63 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3129, 3 => 1088, 4 => -1),
    64 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5238, 3 => 4440, 4 => -1),
    65 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5722, 3 => 4280, 4 => -1),
    66 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3540, 3 => 375, 4 => -1),
    67 => integer_vector_t'(0 => 3, 1 => 13, 2 => 191, 3 => 2782, 4 => -1),
    68 => integer_vector_t'(0 => 3, 1 => 14, 2 => 906, 3 => 4432, 4 => -1),
    69 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3225, 3 => 1111, 4 => -1),
    70 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6296, 3 => 2583, 4 => -1),
    71 => integer_vector_t'(0 => 3, 1 => 17, 2 => 1457, 3 => 903, 4 => -1),
    72 => integer_vector_t'(0 => 3, 1 => 0, 2 => 855, 3 => 4475, 4 => -1),
    73 => integer_vector_t'(0 => 3, 1 => 1, 2 => 4097, 3 => 3970, 4 => -1),
    74 => integer_vector_t'(0 => 3, 1 => 2, 2 => 4433, 3 => 4361, 4 => -1),
    75 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5198, 3 => 541, 4 => -1),
    76 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1146, 3 => 4426, 4 => -1),
    77 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3202, 3 => 2902, 4 => -1),
    78 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2724, 3 => 525, 4 => -1),
    79 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1083, 3 => 4124, 4 => -1),
    80 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2326, 3 => 6003, 4 => -1),
    81 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5605, 3 => 5990, 4 => -1),
    82 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4376, 3 => 1579, 4 => -1),
    83 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4407, 3 => 984, 4 => -1),
    84 => integer_vector_t'(0 => 3, 1 => 12, 2 => 1332, 3 => 6163, 4 => -1),
    85 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5359, 3 => 3975, 4 => -1),
    86 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1907, 3 => 1854, 4 => -1),
    87 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3601, 3 => 5748, 4 => -1),
    88 => integer_vector_t'(0 => 3, 1 => 16, 2 => 6056, 3 => 3266, 4 => -1),
    89 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3322, 3 => 4085, 4 => -1),
    90 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1768, 3 => 3244, 4 => -1),
    91 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2149, 3 => 144, 4 => -1),
    92 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1589, 3 => 4291, 4 => -1),
    93 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5154, 3 => 1252, 4 => -1),
    94 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1855, 3 => 5939, 4 => -1),
    95 => integer_vector_t'(0 => 3, 1 => 5, 2 => 4820, 3 => 2706, 4 => -1),
    96 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1475, 3 => 3360, 4 => -1),
    97 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4266, 3 => 693, 4 => -1),
    98 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4156, 3 => 2018, 4 => -1),
    99 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2103, 3 => 752, 4 => -1),
    100 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3710, 3 => 3853, 4 => -1),
    101 => integer_vector_t'(0 => 3, 1 => 11, 2 => 5123, 3 => 931, 4 => -1),
    102 => integer_vector_t'(0 => 3, 1 => 12, 2 => 6146, 3 => 3323, 4 => -1),
    103 => integer_vector_t'(0 => 3, 1 => 13, 2 => 1939, 3 => 5002, 4 => -1),
    104 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5140, 3 => 1437, 4 => -1),
    105 => integer_vector_t'(0 => 3, 1 => 15, 2 => 1263, 3 => 293, 4 => -1),
    106 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5949, 3 => 4665, 4 => -1),
    107 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4548, 3 => 6380, 4 => -1),
    108 => integer_vector_t'(0 => 3, 1 => 0, 2 => 3171, 3 => 4690, 4 => -1),
    109 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5204, 3 => 2114, 4 => -1),
    110 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6384, 3 => 5565, 4 => -1),
    111 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5722, 3 => 1757, 4 => -1),
    112 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2805, 3 => 6264, 4 => -1),
    113 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1202, 3 => 2616, 4 => -1),
    114 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1018, 3 => 3244, 4 => -1),
    115 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4018, 3 => 5289, 4 => -1),
    116 => integer_vector_t'(0 => 3, 1 => 8, 2 => 2257, 3 => 3067, 4 => -1),
    117 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2483, 3 => 3073, 4 => -1),
    118 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1196, 3 => 5329, 4 => -1),
    119 => integer_vector_t'(0 => 3, 1 => 11, 2 => 649, 3 => 3918, 4 => -1),
    120 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3791, 3 => 4581, 4 => -1),
    121 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5028, 3 => 3803, 4 => -1),
    122 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3119, 3 => 3506, 4 => -1),
    123 => integer_vector_t'(0 => 3, 1 => 15, 2 => 4779, 3 => 431, 4 => -1),
    124 => integer_vector_t'(0 => 3, 1 => 16, 2 => 3888, 3 => 5510, 4 => -1),
    125 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4387, 3 => 4084, 4 => -1),
    126 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5836, 3 => 1692, 4 => -1),
    127 => integer_vector_t'(0 => 3, 1 => 1, 2 => 5126, 3 => 1078, 4 => -1),
    128 => integer_vector_t'(0 => 3, 1 => 2, 2 => 5721, 3 => 6165, 4 => -1),
    129 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3540, 3 => 2499, 4 => -1),
    130 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2225, 3 => 6348, 4 => -1),
    131 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1044, 3 => 1484, 4 => -1),
    132 => integer_vector_t'(0 => 3, 1 => 6, 2 => 6323, 3 => 4042, 4 => -1),
    133 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1313, 3 => 5603, 4 => -1),
    134 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1303, 3 => 3496, 4 => -1),
    135 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3516, 3 => 3639, 4 => -1),
    136 => integer_vector_t'(0 => 3, 1 => 10, 2 => 5161, 3 => 2293, 4 => -1),
    137 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4682, 3 => 3845, 4 => -1),
    138 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3045, 3 => 643, 4 => -1),
    139 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2818, 3 => 2616, 4 => -1),
    140 => integer_vector_t'(0 => 3, 1 => 14, 2 => 3267, 3 => 649, 4 => -1),
    141 => integer_vector_t'(0 => 3, 1 => 15, 2 => 6236, 3 => 593, 4 => -1),
    142 => integer_vector_t'(0 => 3, 1 => 16, 2 => 646, 3 => 2948, 4 => -1),
    143 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4213, 3 => 1442, 4 => -1),
    144 => integer_vector_t'(0 => 3, 1 => 0, 2 => 5779, 3 => 1596, 4 => -1),
    145 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2403, 3 => 1237, 4 => -1),
    146 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2217, 3 => 1514, 4 => -1),
    147 => integer_vector_t'(0 => 3, 1 => 3, 2 => 5609, 3 => 716, 4 => -1),
    148 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5155, 3 => 3858, 4 => -1),
    149 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1517, 3 => 1312, 4 => -1),
    150 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2554, 3 => 3158, 4 => -1),
    151 => integer_vector_t'(0 => 3, 1 => 7, 2 => 5280, 3 => 2643, 4 => -1),
    152 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4990, 3 => 1353, 4 => -1),
    153 => integer_vector_t'(0 => 3, 1 => 9, 2 => 5648, 3 => 1170, 4 => -1),
    154 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1152, 3 => 4366, 4 => -1),
    155 => integer_vector_t'(0 => 3, 1 => 11, 2 => 3561, 3 => 5368, 4 => -1),
    156 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3581, 3 => 1411, 4 => -1),
    157 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5647, 3 => 4661, 4 => -1),
    158 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1542, 3 => 5401, 4 => -1),
    159 => integer_vector_t'(0 => 3, 1 => 15, 2 => 5078, 3 => 2687, 4 => -1),
    160 => integer_vector_t'(0 => 3, 1 => 16, 2 => 316, 3 => 1755, 4 => -1),
    161 => integer_vector_t'(0 => 3, 1 => 17, 2 => 3392, 3 => 1991, 4 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_2.csv, table is 20x100 (250.0 bytes)
  -- Resource estimation: 6 x 18 kB BRAMs or 3 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_2_COLUMN_WIDTHS : integer_vector_t := (0 => 3, 1 => 5, 2 => 14, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_2 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 19)(0 to 8)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 8, 1 => 20, 2 => 712, 3 => 2386, 4 => 6354, 5 => 4061, 6 => 1062, 7 => 5045, 8 => 5158),
    1 => integer_vector_t'(0 => 8, 1 => 21, 2 => 2543, 3 => 5748, 4 => 4822, 5 => 2348, 6 => 3089, 7 => 6328, 8 => 5876),
    2 => integer_vector_t'(0 => 8, 1 => 22, 2 => 926, 3 => 5701, 4 => 269, 5 => 3693, 6 => 2438, 7 => 3190, 8 => 3507),
    3 => integer_vector_t'(0 => 8, 1 => 23, 2 => 2802, 3 => 4520, 4 => 3577, 5 => 5324, 6 => 1091, 7 => 4667, 8 => 4449),
    4 => integer_vector_t'(0 => 8, 1 => 24, 2 => 5140, 3 => 2003, 4 => 1263, 5 => 4742, 6 => 6497, 7 => 1185, 8 => 6202),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 4046, 3 => 6934, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2855, 3 => 66, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 6694, 3 => 212, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3439, 3 => 1158, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 3850, 3 => 4422, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 5924, 3 => 290, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 1467, 3 => 4049, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 7820, 3 => 2242, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4606, 3 => 3080, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4633, 3 => 7877, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3884, 3 => 6868, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 11, 2 => 8935, 3 => 4996, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3028, 3 => 764, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 13, 2 => 5988, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 14, 2 => 7411, 3 => 3450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_3.csv, table is 15x170 (318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 13, 9 => 14, 10 => 14, 11 => 14, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_3 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 14)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 416, 2 => 8909, 3 => 4156, 4 => 3216, 5 => 3112, 6 => 2560, 7 => 2912, 8 => 6405, 9 => 8593, 10 => 4969, 11 => 6723, 12 => 6912),
    1 => integer_vector_t'(0 => 12, 1 => 8978, 2 => 3011, 3 => 4339, 4 => 9312, 5 => 6396, 6 => 2957, 7 => 7288, 8 => 5485, 9 => 6031, 10 => 10218, 11 => 2226, 12 => 3575),
    2 => integer_vector_t'(0 => 12, 1 => 3383, 2 => 10059, 3 => 1114, 4 => 10008, 5 => 10147, 6 => 9384, 7 => 4290, 8 => 434, 9 => 5139, 10 => 3536, 11 => 1965, 12 => 2291),
    3 => integer_vector_t'(0 => 12, 1 => 2797, 2 => 3693, 3 => 7615, 4 => 7077, 5 => 743, 6 => 1941, 7 => 8716, 8 => 6215, 9 => 3840, 10 => 5140, 11 => 4582, 12 => 5420),
    4 => integer_vector_t'(0 => 12, 1 => 6110, 2 => 8551, 3 => 1515, 4 => 7404, 5 => 4879, 6 => 4946, 7 => 5383, 8 => 1831, 9 => 3441, 10 => 9569, 11 => 10472, 12 => 4306),
    5 => integer_vector_t'(0 => 3, 1 => 1505, 2 => 5682, 3 => 7778, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 7172, 2 => 6830, 3 => 6623, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7281, 2 => 3941, 3 => 3505, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 10270, 2 => 8669, 3 => 914, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 3622, 2 => 7563, 3 => 9388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 9930, 2 => 5058, 3 => 4554, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 4844, 2 => 9609, 3 => 2707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 6883, 2 => 3237, 3 => 1714, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4768, 2 => 3878, 3 => 10017, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 10127, 2 => 3334, 3 => 8267, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C1_4.csv, table is 9x171 (192.375 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C1_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 13, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C1_4 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 8)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 6295, 2 => 9626, 3 => 304, 4 => 7695, 5 => 4839, 6 => 4936, 7 => 1660, 8 => 144, 9 => 11203, 10 => 5567, 11 => 6347, 12 => 12557),
    1 => integer_vector_t'(0 => 12, 1 => 10691, 2 => 4988, 3 => 3859, 4 => 3734, 5 => 3071, 6 => 3494, 7 => 7687, 8 => 10313, 9 => 5964, 10 => 8069, 11 => 8296, 12 => 11090),
    2 => integer_vector_t'(0 => 12, 1 => 10774, 2 => 3613, 3 => 5208, 4 => 11177, 5 => 7676, 6 => 3549, 7 => 8746, 8 => 6583, 9 => 7239, 10 => 12265, 11 => 2674, 12 => 4292),
    3 => integer_vector_t'(0 => 12, 1 => 11869, 2 => 3708, 3 => 5981, 4 => 8718, 5 => 4908, 6 => 10650, 7 => 6805, 8 => 3334, 9 => 2627, 10 => 10461, 11 => 9285, 12 => 11120),
    4 => integer_vector_t'(0 => 3, 1 => 7844, 2 => 3079, 3 => 10773, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 3385, 2 => 10854, 3 => 5747, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1360, 2 => 12010, 3 => 12202, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 6189, 2 => 4241, 3 => 2343, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9840, 2 => 12726, 3 => 4977, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_3.csv, table is 30x156 (585.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_3_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 13, 4 => 12, 5 => 12, 6 => 11, 7 => 12, 8 => 13, 9 => 12, 10 => 13, 11 => 12, 12 => 13, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_3 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 29)(0 to 13)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 13, 1 => 0, 2 => 2084, 3 => 1613, 4 => 1548, 5 => 1286, 6 => 1460, 7 => 3196, 8 => 4297, 9 => 2481, 10 => 3369, 11 => 3451, 12 => 4620, 13 => 2622),
    1 => integer_vector_t'(0 => 13, 1 => 1, 2 => 122, 3 => 1516, 4 => 3448, 5 => 2880, 6 => 1407, 7 => 1847, 8 => 3799, 9 => 3529, 10 => 373, 11 => 971, 12 => 4358, 13 => 3108),
    2 => integer_vector_t'(0 => 13, 1 => 2, 2 => 259, 3 => 3399, 4 => 929, 5 => 2650, 6 => 864, 7 => 3996, 8 => 3833, 9 => 107, 10 => 5287, 11 => 164, 12 => 3125, 13 => 2350),
    3 => integer_vector_t'(0 => 3, 1 => 3, 2 => 342, 3 => 3529, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 4, 2 => 4198, 3 => 2147, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1880, 3 => 4836, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3864, 3 => 4910, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 7, 2 => 243, 3 => 1542, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3011, 3 => 1436, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2167, 3 => 2512, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4606, 3 => 1003, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2835, 3 => 705, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3426, 3 => 2365, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 13, 2 => 3848, 3 => 2474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1360, 3 => 1743, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 163, 3 => 2536, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2583, 3 => 1180, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1542, 3 => 509, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 4418, 3 => 1005, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5212, 3 => 5117, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2155, 3 => 2922, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 347, 3 => 2696, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 226, 3 => 4296, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1560, 3 => 487, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3926, 3 => 1640, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 10, 2 => 149, 3 => 2928, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2364, 3 => 563, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 12, 2 => 635, 3 => 688, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 13, 2 => 231, 3 => 1684, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 14, 2 => 1129, 3 => 3894, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C2_5.csv, table is 18x168 (378.0 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C2_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 13, 8 => 13, 9 => 13, 10 => 14, 11 => 13, 12 => 14);

  constant LDPC_TABLE_FECFRAME_SHORT_C2_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 17)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 5650, 2 => 4143, 3 => 8750, 4 => 583, 5 => 6720, 6 => 8071, 7 => 635, 8 => 1767, 9 => 1344, 10 => 6922, 11 => 738, 12 => 6658),
    1 => integer_vector_t'(0 => 12, 1 => 5696, 2 => 1685, 3 => 3207, 4 => 415, 5 => 7019, 6 => 5023, 7 => 5608, 8 => 2605, 9 => 857, 10 => 6915, 11 => 1770, 12 => 8016),
    2 => integer_vector_t'(0 => 12, 1 => 3992, 2 => 771, 3 => 2190, 4 => 7258, 5 => 8970, 6 => 7792, 7 => 1802, 8 => 1866, 9 => 6137, 10 => 8841, 11 => 886, 12 => 1931),
    3 => integer_vector_t'(0 => 12, 1 => 4108, 2 => 3781, 3 => 7577, 4 => 6810, 5 => 9322, 6 => 8226, 7 => 5396, 8 => 5867, 9 => 4428, 10 => 8827, 11 => 7766, 12 => 2254),
    4 => integer_vector_t'(0 => 12, 1 => 4247, 2 => 888, 3 => 4367, 4 => 8821, 5 => 9660, 6 => 324, 7 => 5864, 8 => 4774, 9 => 227, 10 => 7889, 11 => 6405, 12 => 8963),
    5 => integer_vector_t'(0 => 12, 1 => 9693, 2 => 500, 3 => 2520, 4 => 2227, 5 => 1811, 6 => 9330, 7 => 1928, 8 => 5140, 9 => 4030, 10 => 4824, 11 => 806, 12 => 3134),
    6 => integer_vector_t'(0 => 3, 1 => 1652, 2 => 8171, 3 => 1435, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 3366, 2 => 6543, 3 => 3745, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 9286, 2 => 8509, 3 => 4645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 7397, 2 => 5790, 3 => 8972, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 6597, 2 => 4422, 3 => 1799, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 9276, 2 => 4041, 3 => 3847, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 8683, 2 => 7378, 3 => 4946, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 5348, 2 => 1993, 3 => 9186, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 6724, 2 => 9015, 3 => 5646, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 4502, 2 => 4439, 3 => 8474, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 5107, 2 => 7342, 3 => 9442, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 1387, 2 => 8910, 3 => 2660, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_4.csv, table is 33x133 (548.625 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_4_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 4, 2 => 13, 3 => 12, 4 => 13, 5 => 11, 6 => 10, 7 => 12, 8 => 11, 9 => 12, 10 => 10, 11 => 10, 12 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_4 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 32)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 3, 2 => 3198, 3 => 478, 4 => 4207, 5 => 1481, 6 => 1009, 7 => 2616, 8 => 1924, 9 => 3437, 10 => 554, 11 => 683, 12 => 1801),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2681, 3 => 2135, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3107, 3 => 4027, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2637, 3 => 3373, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 3830, 3 => 3449, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 8, 2 => 4129, 3 => 2060, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 9, 2 => 4184, 3 => 2742, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 10, 2 => 3946, 3 => 1070, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 11, 2 => 2239, 3 => 984, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1458, 3 => 3031, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3003, 3 => 1328, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1137, 3 => 1716, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 132, 3 => 3725, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1817, 3 => 638, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1774, 3 => 3447, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3632, 3 => 1257, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 542, 3 => 3694, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1015, 3 => 1945, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 1948, 3 => 412, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 995, 3 => 2238, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4141, 3 => 1907, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2480, 3 => 3079, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 3021, 3 => 1088, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 713, 3 => 1379, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 997, 3 => 3903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2323, 3 => 3361, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1110, 3 => 986, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2532, 3 => 142, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 1690, 3 => 2405, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1298, 3 => 1881, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 9, 2 => 615, 3 => 174, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 10, 2 => 1648, 3 => 3112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 11, 2 => 1415, 3 => 2808, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C3_5.csv, table is 27x160 (540.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C3_5_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 13, 2 => 13, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13, 9 => 13, 10 => 13, 11 => 13, 12 => 13);

  constant LDPC_TABLE_FECFRAME_SHORT_C3_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 26)(0 to 12)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 12, 1 => 2765, 2 => 5713, 3 => 6426, 4 => 3596, 5 => 1374, 6 => 4811, 7 => 2182, 8 => 544, 9 => 3394, 10 => 2840, 11 => 4310, 12 => 771),
    1 => integer_vector_t'(0 => 12, 1 => 4951, 2 => 211, 3 => 2208, 4 => 723, 5 => 1246, 6 => 2928, 7 => 398, 8 => 5739, 9 => 265, 10 => 5601, 11 => 5993, 12 => 2615),
    2 => integer_vector_t'(0 => 12, 1 => 210, 2 => 4730, 3 => 5777, 4 => 3096, 5 => 4282, 6 => 6238, 7 => 4939, 8 => 1119, 9 => 6463, 10 => 5298, 11 => 6320, 12 => 4016),
    3 => integer_vector_t'(0 => 12, 1 => 4167, 2 => 2063, 3 => 4757, 4 => 3157, 5 => 5664, 6 => 3956, 7 => 6045, 8 => 563, 9 => 4284, 10 => 2441, 11 => 3412, 12 => 6334),
    4 => integer_vector_t'(0 => 12, 1 => 4201, 2 => 2428, 3 => 4474, 4 => 59, 5 => 1721, 6 => 736, 7 => 2997, 8 => 428, 9 => 3807, 10 => 1513, 11 => 4732, 12 => 6195),
    5 => integer_vector_t'(0 => 12, 1 => 2670, 2 => 3081, 3 => 5139, 4 => 3736, 5 => 1999, 6 => 5889, 7 => 4362, 8 => 3806, 9 => 4534, 10 => 5409, 11 => 6384, 12 => 5809),
    6 => integer_vector_t'(0 => 12, 1 => 5516, 2 => 1622, 3 => 2906, 4 => 3285, 5 => 1257, 6 => 5797, 7 => 3816, 8 => 817, 9 => 875, 10 => 2311, 11 => 3543, 12 => 1205),
    7 => integer_vector_t'(0 => 12, 1 => 4244, 2 => 2184, 3 => 5415, 4 => 1705, 5 => 5642, 6 => 4886, 7 => 2333, 8 => 287, 9 => 1848, 10 => 1121, 11 => 3595, 12 => 6022),
    8 => integer_vector_t'(0 => 12, 1 => 2142, 2 => 2830, 3 => 4069, 4 => 5654, 5 => 1295, 6 => 2951, 7 => 3919, 8 => 1356, 9 => 884, 10 => 1786, 11 => 396, 12 => 4738),
    9 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2161, 3 => 2653, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1380, 3 => 1461, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2502, 3 => 3707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3971, 3 => 1057, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 4, 2 => 5985, 3 => 6062, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1733, 3 => 6028, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3786, 3 => 1936, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 7, 2 => 4292, 3 => 956, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 8, 2 => 5692, 3 => 3417, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 9, 2 => 266, 3 => 4878, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 10, 2 => 4913, 3 => 3247, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 11, 2 => 4763, 3 => 3937, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 12, 2 => 3590, 3 => 2903, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 13, 2 => 2566, 3 => 4215, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 14, 2 => 5208, 3 => 4707, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 15, 2 => 3940, 3 => 3388, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 16, 2 => 5109, 3 => 4556, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 17, 2 => 4908, 3 => 4177, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C4_5.csv, table is 35x30 (131.25 bytes)
  -- Resource estimation: 2 x 18 kB BRAMs or 1 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C4_5_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 4, 2 => 12, 3 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C4_5 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 34)(0 to 3)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 3, 1 => 5, 2 => 896, 3 => 1565),
    1 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2493, 3 => 184),
    2 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 3210),
    3 => integer_vector_t'(0 => 3, 1 => 8, 2 => 727, 3 => 1339),
    4 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3428, 3 => 612),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2663, 3 => 1947),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 230, 3 => 2695),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2025, 3 => 2794),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3039, 3 => 283),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 862, 3 => 2889),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 376, 3 => 2110),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2034, 3 => 2286),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 951, 3 => 2068),
    13 => integer_vector_t'(0 => 3, 1 => 8, 2 => 3108, 3 => 3542),
    14 => integer_vector_t'(0 => 3, 1 => 9, 2 => 307, 3 => 1421),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2272, 3 => 1197),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1800, 3 => 3280),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 331, 3 => 2308),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 465, 3 => 2552),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1038, 3 => 2479),
    20 => integer_vector_t'(0 => 3, 1 => 5, 2 => 1383, 3 => 343),
    21 => integer_vector_t'(0 => 3, 1 => 6, 2 => 94, 3 => 236),
    22 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2619, 3 => 121),
    23 => integer_vector_t'(0 => 3, 1 => 8, 2 => 1497, 3 => 2774),
    24 => integer_vector_t'(0 => 3, 1 => 9, 2 => 2116, 3 => 1855),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 722, 3 => 1584),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2767, 3 => 1881),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 2701, 3 => 1610),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 3283, 3 => 1732),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 168, 3 => 1099),
    30 => integer_vector_t'(0 => 3, 1 => 5, 2 => 3074, 3 => 243),
    31 => integer_vector_t'(0 => 3, 1 => 6, 2 => 3460, 3 => 945),
    32 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2049, 3 => 1746),
    33 => integer_vector_t'(0 => 3, 1 => 8, 2 => 566, 3 => 1427),
    34 => integer_vector_t'(0 => 3, 1 => 9, 2 => 3545, 3 => 1168)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C5_6.csv, table is 37x139 (642.875 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C5_6_COLUMN_WIDTHS : integer_vector_t := (0 => 4, 1 => 3, 2 => 12, 3 => 12, 4 => 11, 5 => 10, 6 => 10, 7 => 10, 8 => 11, 9 => 9, 10 => 12, 11 => 12, 12 => 11, 13 => 12);

  constant LDPC_TABLE_FECFRAME_SHORT_C5_6 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 36)(0 to 13)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 13, 1 => 3, 2 => 2409, 3 => 499, 4 => 1481, 5 => 908, 6 => 559, 7 => 716, 8 => 1270, 9 => 333, 10 => 2508, 11 => 2264, 12 => 1702, 13 => 2805),
    1 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2447, 3 => 1926, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    2 => integer_vector_t'(0 => 3, 1 => 5, 2 => 414, 3 => 1224, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    3 => integer_vector_t'(0 => 3, 1 => 6, 2 => 2114, 3 => 842, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    4 => integer_vector_t'(0 => 3, 1 => 7, 2 => 212, 3 => 573, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2383, 3 => 2112, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 2286, 3 => 2348, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 545, 3 => 819, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1264, 3 => 143, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1701, 3 => 2258, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 5, 2 => 964, 3 => 166, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 6, 2 => 114, 3 => 2413, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2243, 3 => 81, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1245, 3 => 1581, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 1, 2 => 775, 3 => 169, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1696, 3 => 1104, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1914, 3 => 2831, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 4, 2 => 532, 3 => 1450, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 5, 2 => 91, 3 => 974, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 6, 2 => 497, 3 => 2228, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2326, 3 => 1579, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 0, 2 => 2482, 3 => 256, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1117, 3 => 1261, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1257, 3 => 1658, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1478, 3 => 1225, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 4, 2 => 2511, 3 => 980, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2320, 3 => 2675, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 6, 2 => 435, 3 => 1278, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 7, 2 => 228, 3 => 503, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1885, 3 => 2369, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 1, 2 => 57, 3 => 483, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 2, 2 => 838, 3 => 1050, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1231, 3 => 1990, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1738, 3 => 68, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 5, 2 => 2392, 3 => 951, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 6, 2 => 163, 3 => 645, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 7, 2 => 2644, 3 => 1704, 4 => -1, 5 => -1, 6 => -1, 7 => -1, 8 => -1, 9 => -1, 10 => -1, 11 => -1, 12 => -1, 13 => -1)
  );

  -- From ldpc/ldpc_table_FECFRAME_SHORT_C8_9.csv, table is 40x37 (185.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  constant LDPC_TABLE_FECFRAME_SHORT_C8_9_COLUMN_WIDTHS : integer_vector_t := (0 => 2, 1 => 2, 2 => 11, 3 => 11, 4 => 11);

  constant LDPC_TABLE_FECFRAME_SHORT_C8_9 : integer_2d_array_t
  -- xilinx translate_off
  (0 to 39)(0 to 4)
  -- xilinx translate_on
  := (
    0 => integer_vector_t'(0 => 4, 1 => 0, 2 => 1558, 3 => 712, 4 => 805),
    1 => integer_vector_t'(0 => 4, 1 => 1, 2 => 1450, 3 => 873, 4 => 1337),
    2 => integer_vector_t'(0 => 4, 1 => 2, 2 => 1741, 3 => 1129, 4 => 1184),
    3 => integer_vector_t'(0 => 4, 1 => 3, 2 => 294, 3 => 806, 4 => 1566),
    4 => integer_vector_t'(0 => 4, 1 => 4, 2 => 482, 3 => 605, 4 => 923),
    5 => integer_vector_t'(0 => 3, 1 => 0, 2 => 926, 3 => 1578, 4 => -1),
    6 => integer_vector_t'(0 => 3, 1 => 1, 2 => 777, 3 => 1374, 4 => -1),
    7 => integer_vector_t'(0 => 3, 1 => 2, 2 => 608, 3 => 151, 4 => -1),
    8 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1195, 3 => 210, 4 => -1),
    9 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1484, 3 => 692, 4 => -1),
    10 => integer_vector_t'(0 => 3, 1 => 0, 2 => 427, 3 => 488, 4 => -1),
    11 => integer_vector_t'(0 => 3, 1 => 1, 2 => 828, 3 => 1124, 4 => -1),
    12 => integer_vector_t'(0 => 3, 1 => 2, 2 => 874, 3 => 1366, 4 => -1),
    13 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1500, 3 => 835, 4 => -1),
    14 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1496, 3 => 502, 4 => -1),
    15 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1006, 3 => 1701, 4 => -1),
    16 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1155, 3 => 97, 4 => -1),
    17 => integer_vector_t'(0 => 3, 1 => 2, 2 => 657, 3 => 1403, 4 => -1),
    18 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1453, 3 => 624, 4 => -1),
    19 => integer_vector_t'(0 => 3, 1 => 4, 2 => 429, 3 => 1495, 4 => -1),
    20 => integer_vector_t'(0 => 3, 1 => 0, 2 => 809, 3 => 385, 4 => -1),
    21 => integer_vector_t'(0 => 3, 1 => 1, 2 => 367, 3 => 151, 4 => -1),
    22 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1323, 3 => 202, 4 => -1),
    23 => integer_vector_t'(0 => 3, 1 => 3, 2 => 960, 3 => 318, 4 => -1),
    24 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1451, 3 => 1039, 4 => -1),
    25 => integer_vector_t'(0 => 3, 1 => 0, 2 => 1098, 3 => 1722, 4 => -1),
    26 => integer_vector_t'(0 => 3, 1 => 1, 2 => 1015, 3 => 1428, 4 => -1),
    27 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1261, 3 => 1564, 4 => -1),
    28 => integer_vector_t'(0 => 3, 1 => 3, 2 => 544, 3 => 1190, 4 => -1),
    29 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1472, 3 => 1246, 4 => -1),
    30 => integer_vector_t'(0 => 3, 1 => 0, 2 => 508, 3 => 630, 4 => -1),
    31 => integer_vector_t'(0 => 3, 1 => 1, 2 => 421, 3 => 1704, 4 => -1),
    32 => integer_vector_t'(0 => 3, 1 => 2, 2 => 284, 3 => 898, 4 => -1),
    33 => integer_vector_t'(0 => 3, 1 => 3, 2 => 392, 3 => 577, 4 => -1),
    34 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1155, 3 => 556, 4 => -1),
    35 => integer_vector_t'(0 => 3, 1 => 0, 2 => 631, 3 => 1000, 4 => -1),
    36 => integer_vector_t'(0 => 3, 1 => 1, 2 => 732, 3 => 1368, 4 => -1),
    37 => integer_vector_t'(0 => 3, 1 => 2, 2 => 1328, 3 => 329, 4 => -1),
    38 => integer_vector_t'(0 => 3, 1 => 3, 2 => 1515, 3 => 506, 4 => -1),
    39 => integer_vector_t'(0 => 3, 1 => 4, 2 => 1104, 3 => 1172, 4 => -1)
  );


end package ldpc_tables_pkg;